// Benchmark "miter" written by ABC on Wed Apr 26 17:16:06 2017

module miter ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    po0  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19;
  output po0;
  wire n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
    n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
    n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
    n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
    n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011;
  assign n22 = pi16 & pi17;
  assign n23 = pi14 & pi19;
  assign n24 = n22 & n23;
  assign n25 = pi17 & pi18;
  assign n26 = ~n24 & n25;
  assign n27 = n24 & ~n25;
  assign n28 = ~n26 & ~n27;
  assign n29 = pi16 & pi19;
  assign n30 = ~n28 & n29;
  assign n31 = pi18 & pi19;
  assign n32 = n30 & ~n31;
  assign n33 = ~n30 & n31;
  assign n34 = ~n32 & ~n33;
  assign n35 = n24 & n25;
  assign n36 = ~n34 & ~n35;
  assign n37 = n34 & n35;
  assign n38 = ~n36 & ~n37;
  assign n39 = pi15 & pi16;
  assign n40 = pi12 & pi19;
  assign n41 = n39 & n40;
  assign n42 = pi14 & pi17;
  assign n43 = n40 & n42;
  assign n44 = ~n41 & ~n43;
  assign n45 = n39 & n42;
  assign n46 = n44 & ~n45;
  assign n47 = pi15 & pi18;
  assign n48 = n46 & n47;
  assign n49 = ~n46 & ~n47;
  assign n50 = ~n48 & ~n49;
  assign n51 = n22 & ~n23;
  assign n52 = ~n22 & n23;
  assign n53 = ~n51 & ~n52;
  assign n54 = ~n50 & ~n53;
  assign n55 = ~n46 & n47;
  assign n56 = n54 & n55;
  assign n57 = ~n28 & ~n29;
  assign n58 = n28 & n29;
  assign n59 = ~n57 & ~n58;
  assign n60 = n55 & ~n59;
  assign n61 = ~n56 & ~n60;
  assign n62 = n54 & ~n59;
  assign n63 = n61 & ~n62;
  assign n64 = n38 & n63;
  assign n65 = n54 & n59;
  assign n66 = ~n54 & ~n59;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~n55 & ~n67;
  assign n69 = n55 & n67;
  assign n70 = ~n68 & ~n69;
  assign n71 = pi13 & pi16;
  assign n72 = pi12 & pi17;
  assign n73 = n71 & n72;
  assign n74 = pi14 & pi15;
  assign n75 = n72 & n74;
  assign n76 = ~n73 & ~n75;
  assign n77 = n71 & n74;
  assign n78 = n76 & ~n77;
  assign n79 = pi13 & pi18;
  assign n80 = n78 & n79;
  assign n81 = ~n78 & ~n79;
  assign n82 = ~n80 & ~n81;
  assign n83 = n39 & ~n42;
  assign n84 = ~n39 & n42;
  assign n85 = ~n83 & ~n84;
  assign n86 = ~n40 & ~n85;
  assign n87 = n40 & n85;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n82 & ~n88;
  assign n90 = n71 & ~n74;
  assign n91 = ~n71 & n74;
  assign n92 = ~n90 & ~n91;
  assign n93 = ~n72 & ~n92;
  assign n94 = n72 & n92;
  assign n95 = ~n93 & ~n94;
  assign n96 = pi10 & pi19;
  assign n97 = ~n95 & n96;
  assign n98 = pi10 & pi17;
  assign n99 = pi08 & pi19;
  assign n100 = n98 & n99;
  assign n101 = n96 & n100;
  assign n102 = ~n97 & ~n101;
  assign n103 = ~n95 & n100;
  assign n104 = n102 & ~n103;
  assign n105 = ~n88 & ~n104;
  assign n106 = ~n89 & ~n105;
  assign n107 = ~n82 & ~n104;
  assign n108 = n106 & ~n107;
  assign n109 = ~n78 & n79;
  assign n110 = ~n108 & n109;
  assign n111 = ~n50 & n53;
  assign n112 = n50 & ~n53;
  assign n113 = ~n111 & ~n112;
  assign n114 = n109 & ~n113;
  assign n115 = ~n110 & ~n114;
  assign n116 = ~n108 & ~n113;
  assign n117 = n115 & ~n116;
  assign n118 = n70 & n117;
  assign n119 = ~n108 & n113;
  assign n120 = n108 & ~n113;
  assign n121 = ~n119 & ~n120;
  assign n122 = ~n109 & ~n121;
  assign n123 = n109 & n121;
  assign n124 = ~n122 & ~n123;
  assign n125 = pi11 & pi16;
  assign n126 = pi12 & pi15;
  assign n127 = n125 & n126;
  assign n128 = pi13 & pi14;
  assign n129 = n126 & n128;
  assign n130 = ~n127 & ~n129;
  assign n131 = n125 & n128;
  assign n132 = n130 & ~n131;
  assign n133 = pi11 & pi18;
  assign n134 = n132 & n133;
  assign n135 = ~n132 & ~n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = ~n95 & ~n100;
  assign n138 = n95 & n100;
  assign n139 = ~n137 & ~n138;
  assign n140 = ~n96 & ~n139;
  assign n141 = n96 & n139;
  assign n142 = ~n140 & ~n141;
  assign n143 = ~n136 & ~n142;
  assign n144 = n125 & ~n128;
  assign n145 = ~n125 & n128;
  assign n146 = ~n144 & ~n145;
  assign n147 = ~n126 & ~n146;
  assign n148 = n126 & n146;
  assign n149 = ~n147 & ~n148;
  assign n150 = n98 & ~n99;
  assign n151 = ~n98 & n99;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~n149 & ~n152;
  assign n154 = pi10 & pi15;
  assign n155 = pi06 & pi19;
  assign n156 = n154 & n155;
  assign n157 = pi08 & pi17;
  assign n158 = n155 & n157;
  assign n159 = ~n156 & ~n158;
  assign n160 = n154 & n157;
  assign n161 = n159 & ~n160;
  assign n162 = ~n152 & ~n161;
  assign n163 = ~n153 & ~n162;
  assign n164 = ~n149 & ~n161;
  assign n165 = n163 & ~n164;
  assign n166 = ~n142 & ~n165;
  assign n167 = ~n143 & ~n166;
  assign n168 = ~n136 & ~n165;
  assign n169 = n167 & ~n168;
  assign n170 = ~n132 & n133;
  assign n171 = ~n169 & n170;
  assign n172 = ~n82 & n104;
  assign n173 = n82 & ~n104;
  assign n174 = ~n172 & ~n173;
  assign n175 = n88 & ~n174;
  assign n176 = ~n88 & n174;
  assign n177 = ~n175 & ~n176;
  assign n178 = n170 & ~n177;
  assign n179 = ~n171 & ~n178;
  assign n180 = ~n169 & ~n177;
  assign n181 = n179 & ~n180;
  assign n182 = n124 & n181;
  assign n183 = ~n118 & ~n182;
  assign n184 = ~n64 & n183;
  assign n185 = ~n169 & n177;
  assign n186 = n169 & ~n177;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~n170 & ~n187;
  assign n189 = n170 & n187;
  assign n190 = ~n188 & ~n189;
  assign n191 = pi09 & pi16;
  assign n192 = pi12 & pi13;
  assign n193 = n191 & n192;
  assign n194 = pi11 & pi14;
  assign n195 = n192 & n194;
  assign n196 = ~n193 & ~n195;
  assign n197 = n191 & n194;
  assign n198 = n196 & ~n197;
  assign n199 = pi09 & pi18;
  assign n200 = n198 & n199;
  assign n201 = ~n198 & ~n199;
  assign n202 = ~n200 & ~n201;
  assign n203 = ~n149 & n161;
  assign n204 = n149 & ~n161;
  assign n205 = ~n203 & ~n204;
  assign n206 = n152 & ~n205;
  assign n207 = ~n152 & n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n202 & ~n208;
  assign n210 = n191 & ~n194;
  assign n211 = ~n191 & n194;
  assign n212 = ~n210 & ~n211;
  assign n213 = ~n192 & ~n212;
  assign n214 = n192 & n212;
  assign n215 = ~n213 & ~n214;
  assign n216 = n154 & ~n157;
  assign n217 = ~n154 & n157;
  assign n218 = ~n216 & ~n217;
  assign n219 = ~n155 & ~n218;
  assign n220 = n155 & n218;
  assign n221 = ~n219 & ~n220;
  assign n222 = ~n215 & ~n221;
  assign n223 = pi10 & pi13;
  assign n224 = pi06 & pi17;
  assign n225 = n223 & n224;
  assign n226 = pi08 & pi15;
  assign n227 = n224 & n226;
  assign n228 = ~n225 & ~n227;
  assign n229 = n223 & n226;
  assign n230 = n228 & ~n229;
  assign n231 = ~n221 & ~n230;
  assign n232 = ~n222 & ~n231;
  assign n233 = ~n215 & ~n230;
  assign n234 = n232 & ~n233;
  assign n235 = ~n208 & ~n234;
  assign n236 = ~n209 & ~n235;
  assign n237 = ~n202 & ~n234;
  assign n238 = n236 & ~n237;
  assign n239 = ~n198 & n199;
  assign n240 = ~n238 & n239;
  assign n241 = ~n136 & n165;
  assign n242 = n136 & ~n165;
  assign n243 = ~n241 & ~n242;
  assign n244 = n142 & ~n243;
  assign n245 = ~n142 & n243;
  assign n246 = ~n244 & ~n245;
  assign n247 = n239 & ~n246;
  assign n248 = ~n240 & ~n247;
  assign n249 = ~n238 & ~n246;
  assign n250 = n248 & ~n249;
  assign n251 = n190 & n250;
  assign n252 = ~n238 & n246;
  assign n253 = n238 & ~n246;
  assign n254 = ~n252 & ~n253;
  assign n255 = ~n239 & ~n254;
  assign n256 = n239 & n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = pi05 & pi18;
  assign n259 = pi02 & pi19;
  assign n260 = pi04 & pi17;
  assign n261 = n259 & n260;
  assign n262 = n258 & n261;
  assign n263 = pi04 & pi19;
  assign n264 = n258 & n263;
  assign n265 = ~n262 & ~n264;
  assign n266 = n261 & n263;
  assign n267 = n265 & ~n266;
  assign n268 = pi07 & pi18;
  assign n269 = ~n267 & ~n268;
  assign n270 = n267 & n268;
  assign n271 = ~n269 & ~n270;
  assign n272 = pi07 & pi16;
  assign n273 = pi11 & pi12;
  assign n274 = n272 & n273;
  assign n275 = pi09 & pi14;
  assign n276 = n273 & n275;
  assign n277 = ~n274 & ~n276;
  assign n278 = n272 & n275;
  assign n279 = n277 & ~n278;
  assign n280 = ~n271 & n279;
  assign n281 = n271 & ~n279;
  assign n282 = ~n280 & ~n281;
  assign n283 = ~n215 & n230;
  assign n284 = n215 & ~n230;
  assign n285 = ~n283 & ~n284;
  assign n286 = n221 & ~n285;
  assign n287 = ~n221 & n285;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~n282 & ~n288;
  assign n290 = n272 & ~n275;
  assign n291 = ~n272 & n275;
  assign n292 = ~n290 & ~n291;
  assign n293 = ~n273 & ~n292;
  assign n294 = n273 & n292;
  assign n295 = ~n293 & ~n294;
  assign n296 = n223 & ~n226;
  assign n297 = ~n223 & n226;
  assign n298 = ~n296 & ~n297;
  assign n299 = ~n224 & ~n298;
  assign n300 = n224 & n298;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~n295 & ~n301;
  assign n303 = pi10 & pi11;
  assign n304 = pi06 & pi15;
  assign n305 = n303 & n304;
  assign n306 = pi08 & pi13;
  assign n307 = n304 & n306;
  assign n308 = ~n305 & ~n307;
  assign n309 = n303 & n306;
  assign n310 = n308 & ~n309;
  assign n311 = ~n301 & ~n310;
  assign n312 = ~n302 & ~n311;
  assign n313 = ~n295 & ~n310;
  assign n314 = n312 & ~n313;
  assign n315 = ~n288 & ~n314;
  assign n316 = ~n289 & ~n315;
  assign n317 = ~n282 & ~n314;
  assign n318 = n316 & ~n317;
  assign n319 = ~n267 & ~n279;
  assign n320 = n268 & ~n279;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~n267 & n268;
  assign n323 = n321 & ~n322;
  assign n324 = ~n318 & ~n323;
  assign n325 = ~n202 & n234;
  assign n326 = n202 & ~n234;
  assign n327 = ~n325 & ~n326;
  assign n328 = n208 & ~n327;
  assign n329 = ~n208 & n327;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~n323 & ~n330;
  assign n332 = ~n324 & ~n331;
  assign n333 = ~n318 & ~n330;
  assign n334 = n332 & ~n333;
  assign n335 = n257 & n334;
  assign n336 = ~n251 & ~n335;
  assign n337 = ~n318 & n330;
  assign n338 = n318 & ~n330;
  assign n339 = ~n337 & ~n338;
  assign n340 = n323 & ~n339;
  assign n341 = ~n323 & n339;
  assign n342 = ~n340 & ~n341;
  assign n343 = n261 & ~n263;
  assign n344 = ~n261 & n263;
  assign n345 = ~n343 & ~n344;
  assign n346 = ~n258 & ~n345;
  assign n347 = n258 & n345;
  assign n348 = ~n346 & ~n347;
  assign n349 = pi03 & pi18;
  assign n350 = pi00 & pi19;
  assign n351 = pi04 & pi15;
  assign n352 = n350 & n351;
  assign n353 = pi02 & pi17;
  assign n354 = n350 & n353;
  assign n355 = ~n352 & ~n354;
  assign n356 = n351 & n353;
  assign n357 = n355 & ~n356;
  assign n358 = n349 & ~n357;
  assign n359 = ~n259 & n260;
  assign n360 = n259 & ~n260;
  assign n361 = ~n359 & ~n360;
  assign n362 = n349 & ~n361;
  assign n363 = ~n358 & ~n362;
  assign n364 = ~n357 & ~n361;
  assign n365 = n363 & ~n364;
  assign n366 = n348 & ~n365;
  assign n367 = ~n348 & n365;
  assign n368 = ~n366 & ~n367;
  assign n369 = pi05 & pi16;
  assign n370 = pi09 & pi12;
  assign n371 = n369 & n370;
  assign n372 = pi07 & pi14;
  assign n373 = n370 & n372;
  assign n374 = ~n371 & ~n373;
  assign n375 = n369 & n372;
  assign n376 = n374 & ~n375;
  assign n377 = ~n368 & n376;
  assign n378 = n368 & ~n376;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~n295 & n310;
  assign n381 = n295 & ~n310;
  assign n382 = ~n380 & ~n381;
  assign n383 = n301 & ~n382;
  assign n384 = ~n301 & n382;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n379 & ~n385;
  assign n387 = n369 & ~n372;
  assign n388 = ~n369 & n372;
  assign n389 = ~n387 & ~n388;
  assign n390 = ~n370 & ~n389;
  assign n391 = n370 & n389;
  assign n392 = ~n390 & ~n391;
  assign n393 = n303 & ~n306;
  assign n394 = ~n303 & n306;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~n304 & ~n395;
  assign n397 = n304 & n395;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n392 & ~n398;
  assign n400 = pi06 & pi13;
  assign n401 = pi09 & pi10;
  assign n402 = n400 & n401;
  assign n403 = pi08 & pi11;
  assign n404 = n400 & n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = n401 & n403;
  assign n407 = n405 & ~n406;
  assign n408 = ~n398 & ~n407;
  assign n409 = ~n399 & ~n408;
  assign n410 = ~n392 & ~n407;
  assign n411 = n409 & ~n410;
  assign n412 = ~n385 & ~n411;
  assign n413 = ~n386 & ~n412;
  assign n414 = ~n379 & ~n411;
  assign n415 = n413 & ~n414;
  assign n416 = ~n365 & ~n376;
  assign n417 = ~n348 & ~n376;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n348 & ~n365;
  assign n420 = n418 & ~n419;
  assign n421 = ~n415 & ~n420;
  assign n422 = ~n282 & n314;
  assign n423 = n282 & ~n314;
  assign n424 = ~n422 & ~n423;
  assign n425 = n288 & ~n424;
  assign n426 = ~n288 & n424;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~n420 & ~n427;
  assign n429 = ~n421 & ~n428;
  assign n430 = ~n415 & ~n427;
  assign n431 = n429 & ~n430;
  assign n432 = n342 & n431;
  assign n433 = ~n415 & n427;
  assign n434 = n415 & ~n427;
  assign n435 = ~n433 & ~n434;
  assign n436 = n420 & ~n435;
  assign n437 = ~n420 & n435;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n357 & n361;
  assign n440 = n357 & ~n361;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~n349 & ~n441;
  assign n443 = n349 & n441;
  assign n444 = ~n442 & ~n443;
  assign n445 = pi01 & pi18;
  assign n446 = pi00 & pi17;
  assign n447 = pi04 & pi13;
  assign n448 = n446 & n447;
  assign n449 = pi02 & pi15;
  assign n450 = n446 & n449;
  assign n451 = ~n448 & ~n450;
  assign n452 = n447 & n449;
  assign n453 = n451 & ~n452;
  assign n454 = n445 & ~n453;
  assign n455 = n351 & ~n353;
  assign n456 = ~n351 & n353;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~n350 & ~n457;
  assign n459 = n350 & n457;
  assign n460 = ~n458 & ~n459;
  assign n461 = n445 & ~n460;
  assign n462 = ~n454 & ~n461;
  assign n463 = ~n453 & ~n460;
  assign n464 = n462 & ~n463;
  assign n465 = n444 & ~n464;
  assign n466 = ~n444 & n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = pi07 & pi12;
  assign n469 = pi03 & pi16;
  assign n470 = n468 & n469;
  assign n471 = pi05 & pi14;
  assign n472 = n468 & n471;
  assign n473 = ~n470 & ~n472;
  assign n474 = n469 & n471;
  assign n475 = n473 & ~n474;
  assign n476 = ~n467 & n475;
  assign n477 = n467 & ~n475;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~n392 & n407;
  assign n480 = n392 & ~n407;
  assign n481 = ~n479 & ~n480;
  assign n482 = n398 & ~n481;
  assign n483 = ~n398 & n481;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n478 & ~n484;
  assign n486 = n469 & ~n471;
  assign n487 = ~n469 & n471;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~n468 & ~n488;
  assign n490 = n468 & n488;
  assign n491 = ~n489 & ~n490;
  assign n492 = n401 & ~n403;
  assign n493 = ~n401 & n403;
  assign n494 = ~n492 & ~n493;
  assign n495 = ~n400 & ~n494;
  assign n496 = n400 & n494;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n491 & ~n497;
  assign n499 = pi06 & pi11;
  assign n500 = pi07 & pi10;
  assign n501 = n499 & n500;
  assign n502 = pi08 & pi09;
  assign n503 = n499 & n502;
  assign n504 = ~n501 & ~n503;
  assign n505 = n500 & n502;
  assign n506 = n504 & ~n505;
  assign n507 = ~n497 & ~n506;
  assign n508 = ~n498 & ~n507;
  assign n509 = ~n491 & ~n506;
  assign n510 = n508 & ~n509;
  assign n511 = ~n484 & ~n510;
  assign n512 = ~n485 & ~n511;
  assign n513 = ~n478 & ~n510;
  assign n514 = n512 & ~n513;
  assign n515 = ~n464 & ~n475;
  assign n516 = ~n444 & ~n475;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~n444 & ~n464;
  assign n519 = n517 & ~n518;
  assign n520 = ~n514 & ~n519;
  assign n521 = ~n379 & n411;
  assign n522 = n379 & ~n411;
  assign n523 = ~n521 & ~n522;
  assign n524 = n385 & ~n523;
  assign n525 = ~n385 & n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~n519 & ~n526;
  assign n528 = ~n520 & ~n527;
  assign n529 = ~n514 & ~n526;
  assign n530 = n528 & ~n529;
  assign n531 = n438 & n530;
  assign n532 = ~n432 & ~n531;
  assign n533 = n336 & n532;
  assign n534 = ~n514 & n526;
  assign n535 = n514 & ~n526;
  assign n536 = ~n534 & ~n535;
  assign n537 = n519 & ~n536;
  assign n538 = ~n519 & n536;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~n453 & n460;
  assign n541 = n453 & ~n460;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~n445 & ~n542;
  assign n544 = n445 & n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = n447 & ~n449;
  assign n547 = ~n447 & n449;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n446 & ~n548;
  assign n550 = n446 & n548;
  assign n551 = ~n549 & ~n550;
  assign n552 = pi04 & pi11;
  assign n553 = pi00 & pi15;
  assign n554 = n552 & n553;
  assign n555 = pi02 & pi13;
  assign n556 = n553 & n555;
  assign n557 = ~n554 & ~n556;
  assign n558 = n552 & n555;
  assign n559 = n557 & ~n558;
  assign n560 = ~n551 & ~n559;
  assign n561 = n545 & n560;
  assign n562 = ~n545 & ~n560;
  assign n563 = ~n561 & ~n562;
  assign n564 = pi01 & pi16;
  assign n565 = pi05 & pi12;
  assign n566 = n564 & n565;
  assign n567 = pi03 & pi14;
  assign n568 = n565 & n567;
  assign n569 = ~n566 & ~n568;
  assign n570 = n564 & n567;
  assign n571 = n569 & ~n570;
  assign n572 = ~n563 & n571;
  assign n573 = n563 & ~n571;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~n491 & n506;
  assign n576 = n491 & ~n506;
  assign n577 = ~n575 & ~n576;
  assign n578 = n497 & ~n577;
  assign n579 = ~n497 & n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n574 & ~n580;
  assign n582 = n564 & ~n567;
  assign n583 = ~n564 & n567;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n565 & ~n584;
  assign n586 = n565 & n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = n500 & ~n502;
  assign n589 = ~n500 & n502;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n499 & ~n590;
  assign n592 = n499 & n590;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n587 & ~n593;
  assign n595 = pi05 & pi10;
  assign n596 = pi06 & pi09;
  assign n597 = n595 & n596;
  assign n598 = pi07 & pi08;
  assign n599 = n596 & n598;
  assign n600 = ~n597 & ~n599;
  assign n601 = n595 & n598;
  assign n602 = n600 & ~n601;
  assign n603 = ~n593 & ~n602;
  assign n604 = ~n594 & ~n603;
  assign n605 = ~n587 & ~n602;
  assign n606 = n604 & ~n605;
  assign n607 = ~n580 & ~n606;
  assign n608 = ~n581 & ~n607;
  assign n609 = ~n574 & ~n606;
  assign n610 = n608 & ~n609;
  assign n611 = n560 & ~n571;
  assign n612 = ~n545 & ~n571;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n545 & n560;
  assign n615 = n613 & ~n614;
  assign n616 = ~n610 & ~n615;
  assign n617 = ~n478 & n510;
  assign n618 = n478 & ~n510;
  assign n619 = ~n617 & ~n618;
  assign n620 = n484 & ~n619;
  assign n621 = ~n484 & n619;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~n615 & ~n622;
  assign n624 = ~n616 & ~n623;
  assign n625 = ~n610 & ~n622;
  assign n626 = n624 & ~n625;
  assign n627 = n539 & n626;
  assign n628 = ~n610 & n622;
  assign n629 = n610 & ~n622;
  assign n630 = ~n628 & ~n629;
  assign n631 = n615 & ~n630;
  assign n632 = ~n615 & n630;
  assign n633 = ~n631 & ~n632;
  assign n634 = n551 & ~n559;
  assign n635 = ~n551 & n559;
  assign n636 = ~n634 & ~n635;
  assign n637 = pi04 & pi09;
  assign n638 = pi00 & pi13;
  assign n639 = n637 & n638;
  assign n640 = pi02 & pi11;
  assign n641 = n638 & n640;
  assign n642 = ~n639 & ~n641;
  assign n643 = n637 & n640;
  assign n644 = n642 & ~n643;
  assign n645 = n552 & ~n555;
  assign n646 = ~n552 & n555;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n553 & ~n647;
  assign n649 = n553 & n647;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n644 & ~n650;
  assign n652 = n636 & n651;
  assign n653 = ~n636 & ~n651;
  assign n654 = ~n652 & ~n653;
  assign n655 = pi01 & pi14;
  assign n656 = pi03 & pi12;
  assign n657 = n655 & n656;
  assign n658 = ~n654 & ~n657;
  assign n659 = n654 & n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n587 & n602;
  assign n662 = n587 & ~n602;
  assign n663 = ~n661 & ~n662;
  assign n664 = n593 & ~n663;
  assign n665 = ~n593 & n663;
  assign n666 = ~n664 & ~n665;
  assign n667 = ~n660 & ~n666;
  assign n668 = n655 & ~n656;
  assign n669 = ~n655 & n656;
  assign n670 = ~n668 & ~n669;
  assign n671 = n595 & ~n598;
  assign n672 = ~n595 & n598;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~n596 & ~n673;
  assign n675 = n596 & n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n670 & ~n676;
  assign n678 = pi03 & pi10;
  assign n679 = pi06 & pi07;
  assign n680 = n678 & n679;
  assign n681 = pi05 & pi08;
  assign n682 = n679 & n681;
  assign n683 = ~n680 & ~n682;
  assign n684 = n678 & n681;
  assign n685 = n683 & ~n684;
  assign n686 = ~n676 & ~n685;
  assign n687 = ~n677 & ~n686;
  assign n688 = ~n670 & ~n685;
  assign n689 = n687 & ~n688;
  assign n690 = ~n666 & ~n689;
  assign n691 = ~n667 & ~n690;
  assign n692 = ~n660 & ~n689;
  assign n693 = n691 & ~n692;
  assign n694 = n651 & n657;
  assign n695 = ~n636 & n657;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~n636 & n651;
  assign n698 = n696 & ~n697;
  assign n699 = ~n693 & ~n698;
  assign n700 = ~n574 & n606;
  assign n701 = n574 & ~n606;
  assign n702 = ~n700 & ~n701;
  assign n703 = n580 & ~n702;
  assign n704 = ~n580 & n702;
  assign n705 = ~n703 & ~n704;
  assign n706 = ~n698 & ~n705;
  assign n707 = ~n699 & ~n706;
  assign n708 = ~n693 & ~n705;
  assign n709 = n707 & ~n708;
  assign n710 = n633 & n709;
  assign n711 = ~n627 & ~n710;
  assign n712 = ~n693 & n705;
  assign n713 = n693 & ~n705;
  assign n714 = ~n712 & ~n713;
  assign n715 = n698 & ~n714;
  assign n716 = ~n698 & n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = ~n644 & n650;
  assign n719 = n644 & ~n650;
  assign n720 = ~n718 & ~n719;
  assign n721 = pi04 & pi07;
  assign n722 = pi00 & pi11;
  assign n723 = n721 & n722;
  assign n724 = pi02 & pi09;
  assign n725 = n722 & n724;
  assign n726 = ~n723 & ~n725;
  assign n727 = n721 & n724;
  assign n728 = n726 & ~n727;
  assign n729 = n637 & ~n640;
  assign n730 = ~n637 & n640;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~n638 & ~n731;
  assign n733 = n638 & n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n728 & ~n734;
  assign n736 = n720 & n735;
  assign n737 = ~n720 & ~n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~n670 & n685;
  assign n740 = n670 & ~n685;
  assign n741 = ~n739 & ~n740;
  assign n742 = n676 & ~n741;
  assign n743 = ~n676 & n741;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n738 & ~n744;
  assign n746 = n678 & ~n681;
  assign n747 = ~n678 & n681;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n679 & ~n748;
  assign n750 = n679 & n748;
  assign n751 = ~n749 & ~n750;
  assign n752 = pi01 & pi12;
  assign n753 = ~n751 & n752;
  assign n754 = pi01 & pi10;
  assign n755 = pi05 & pi06;
  assign n756 = n754 & n755;
  assign n757 = pi03 & pi08;
  assign n758 = n755 & n757;
  assign n759 = ~n756 & ~n758;
  assign n760 = n754 & n757;
  assign n761 = n759 & ~n760;
  assign n762 = ~n751 & ~n761;
  assign n763 = ~n753 & ~n762;
  assign n764 = n752 & ~n761;
  assign n765 = n763 & ~n764;
  assign n766 = ~n744 & ~n765;
  assign n767 = ~n745 & ~n766;
  assign n768 = ~n738 & ~n765;
  assign n769 = n767 & ~n768;
  assign n770 = ~n720 & n735;
  assign n771 = ~n769 & n770;
  assign n772 = ~n660 & n689;
  assign n773 = n660 & ~n689;
  assign n774 = ~n772 & ~n773;
  assign n775 = n666 & ~n774;
  assign n776 = ~n666 & n774;
  assign n777 = ~n775 & ~n776;
  assign n778 = n770 & ~n777;
  assign n779 = ~n771 & ~n778;
  assign n780 = ~n769 & ~n777;
  assign n781 = n779 & ~n780;
  assign n782 = n717 & n781;
  assign n783 = ~n769 & n777;
  assign n784 = n769 & ~n777;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~n770 & ~n785;
  assign n787 = n770 & n785;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~n728 & n734;
  assign n790 = n728 & ~n734;
  assign n791 = ~n789 & ~n790;
  assign n792 = pi04 & pi05;
  assign n793 = pi00 & pi09;
  assign n794 = n792 & n793;
  assign n795 = pi02 & pi07;
  assign n796 = n793 & n795;
  assign n797 = ~n794 & ~n796;
  assign n798 = n792 & n795;
  assign n799 = n797 & ~n798;
  assign n800 = n721 & ~n724;
  assign n801 = ~n721 & n724;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~n722 & ~n802;
  assign n804 = n722 & n802;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n799 & ~n805;
  assign n807 = n791 & n806;
  assign n808 = ~n791 & ~n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = n752 & n761;
  assign n811 = ~n752 & ~n761;
  assign n812 = ~n810 & ~n811;
  assign n813 = n751 & ~n812;
  assign n814 = ~n751 & n812;
  assign n815 = ~n813 & ~n814;
  assign n816 = ~n809 & ~n815;
  assign n817 = n754 & ~n757;
  assign n818 = ~n754 & n757;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n755 & ~n819;
  assign n821 = n755 & n819;
  assign n822 = ~n820 & ~n821;
  assign n823 = pi01 & pi08;
  assign n824 = pi03 & pi06;
  assign n825 = n823 & n824;
  assign n826 = ~n822 & n825;
  assign n827 = ~n815 & n826;
  assign n828 = ~n816 & ~n827;
  assign n829 = ~n809 & n826;
  assign n830 = n828 & ~n829;
  assign n831 = ~n791 & n806;
  assign n832 = ~n830 & n831;
  assign n833 = ~n738 & n765;
  assign n834 = n738 & ~n765;
  assign n835 = ~n833 & ~n834;
  assign n836 = n744 & ~n835;
  assign n837 = ~n744 & n835;
  assign n838 = ~n836 & ~n837;
  assign n839 = n831 & ~n838;
  assign n840 = ~n832 & ~n839;
  assign n841 = ~n830 & ~n838;
  assign n842 = n840 & ~n841;
  assign n843 = n788 & n842;
  assign n844 = ~n782 & ~n843;
  assign n845 = n711 & n844;
  assign n846 = n533 & n845;
  assign n847 = ~n830 & n838;
  assign n848 = n830 & ~n838;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~n831 & ~n849;
  assign n851 = n831 & n849;
  assign n852 = ~n850 & ~n851;
  assign n853 = ~n799 & n805;
  assign n854 = n799 & ~n805;
  assign n855 = ~n853 & ~n854;
  assign n856 = pi03 & pi04;
  assign n857 = pi00 & pi07;
  assign n858 = n856 & n857;
  assign n859 = pi02 & pi05;
  assign n860 = n857 & n859;
  assign n861 = ~n858 & ~n860;
  assign n862 = n856 & n859;
  assign n863 = n861 & ~n862;
  assign n864 = n792 & ~n795;
  assign n865 = ~n792 & n795;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n793 & ~n866;
  assign n868 = n793 & n866;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~n863 & ~n869;
  assign n871 = n855 & n870;
  assign n872 = ~n855 & ~n870;
  assign n873 = ~n871 & ~n872;
  assign n874 = n822 & n825;
  assign n875 = ~n822 & ~n825;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n873 & ~n876;
  assign n878 = ~n855 & n870;
  assign n879 = n877 & n878;
  assign n880 = ~n809 & ~n826;
  assign n881 = n809 & n826;
  assign n882 = ~n880 & ~n881;
  assign n883 = n815 & ~n882;
  assign n884 = ~n815 & n882;
  assign n885 = ~n883 & ~n884;
  assign n886 = n878 & ~n885;
  assign n887 = ~n879 & ~n886;
  assign n888 = n877 & ~n885;
  assign n889 = n887 & ~n888;
  assign n890 = n852 & n889;
  assign n891 = n877 & n885;
  assign n892 = ~n877 & ~n885;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n878 & ~n893;
  assign n895 = n878 & n893;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~n863 & n869;
  assign n898 = n863 & ~n869;
  assign n899 = ~n897 & ~n898;
  assign n900 = pi01 & pi04;
  assign n901 = pi00 & pi05;
  assign n902 = n900 & n901;
  assign n903 = pi02 & pi03;
  assign n904 = n901 & n903;
  assign n905 = ~n902 & ~n904;
  assign n906 = n900 & n903;
  assign n907 = n905 & ~n906;
  assign n908 = n856 & ~n859;
  assign n909 = ~n856 & n859;
  assign n910 = ~n908 & ~n909;
  assign n911 = ~n857 & ~n910;
  assign n912 = n857 & n910;
  assign n913 = ~n911 & ~n912;
  assign n914 = ~n907 & ~n913;
  assign n915 = n899 & n914;
  assign n916 = ~n899 & ~n914;
  assign n917 = ~n915 & ~n916;
  assign n918 = n823 & ~n824;
  assign n919 = ~n823 & n824;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n917 & ~n920;
  assign n922 = ~n899 & n914;
  assign n923 = n921 & n922;
  assign n924 = ~n873 & n876;
  assign n925 = n873 & ~n876;
  assign n926 = ~n924 & ~n925;
  assign n927 = n922 & ~n926;
  assign n928 = ~n923 & ~n927;
  assign n929 = n921 & ~n926;
  assign n930 = n928 & ~n929;
  assign n931 = n896 & n930;
  assign n932 = ~n890 & ~n931;
  assign n933 = n921 & n926;
  assign n934 = ~n921 & ~n926;
  assign n935 = ~n933 & ~n934;
  assign n936 = ~n922 & ~n935;
  assign n937 = n922 & n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n907 & n913;
  assign n940 = n907 & ~n913;
  assign n941 = ~n939 & ~n940;
  assign n942 = n900 & ~n903;
  assign n943 = ~n900 & n903;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n901 & ~n944;
  assign n946 = n901 & n944;
  assign n947 = ~n945 & ~n946;
  assign n948 = pi00 & pi03;
  assign n949 = pi01 & pi02;
  assign n950 = n948 & n949;
  assign n951 = ~n947 & n950;
  assign n952 = n941 & n951;
  assign n953 = ~n941 & ~n951;
  assign n954 = ~n952 & ~n953;
  assign n955 = pi01 & pi06;
  assign n956 = ~n954 & n955;
  assign n957 = ~n941 & n951;
  assign n958 = n956 & n957;
  assign n959 = ~n917 & n920;
  assign n960 = n917 & ~n920;
  assign n961 = ~n959 & ~n960;
  assign n962 = n957 & ~n961;
  assign n963 = ~n958 & ~n962;
  assign n964 = n956 & ~n961;
  assign n965 = n963 & ~n964;
  assign n966 = ~n938 & ~n965;
  assign n967 = n932 & n966;
  assign n968 = ~n896 & ~n930;
  assign n969 = ~n890 & n968;
  assign n970 = ~n852 & ~n889;
  assign n971 = ~n969 & ~n970;
  assign n972 = ~n967 & n971;
  assign n973 = n846 & ~n972;
  assign n974 = ~n788 & ~n842;
  assign n975 = ~n782 & n974;
  assign n976 = ~n717 & ~n781;
  assign n977 = ~n975 & ~n976;
  assign n978 = n711 & ~n977;
  assign n979 = ~n633 & ~n709;
  assign n980 = ~n627 & n979;
  assign n981 = ~n539 & ~n626;
  assign n982 = ~n980 & ~n981;
  assign n983 = ~n978 & n982;
  assign n984 = n533 & ~n983;
  assign n985 = ~n438 & ~n530;
  assign n986 = ~n432 & n985;
  assign n987 = ~n342 & ~n431;
  assign n988 = ~n986 & ~n987;
  assign n989 = n336 & ~n988;
  assign n990 = ~n257 & ~n334;
  assign n991 = ~n251 & n990;
  assign n992 = ~n190 & ~n250;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n989 & n993;
  assign n995 = ~n984 & n994;
  assign n996 = ~n973 & n995;
  assign n997 = n184 & ~n996;
  assign n998 = ~n124 & ~n181;
  assign n999 = ~n118 & n998;
  assign n1000 = ~n70 & ~n117;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = ~n64 & ~n1001;
  assign n1003 = ~n38 & ~n63;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = ~n997 & n1004;
  assign n1006 = n30 & n35;
  assign n1007 = n31 & n35;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = n30 & n31;
  assign n1010 = n1008 & ~n1009;
  assign n1011 = ~n1005 & n1010;
  assign n1012 = n1005 & ~n1010;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = n224 & n263;
  assign n1015 = ~n266 & ~n1014;
  assign n1016 = n224 & n261;
  assign n1017 = n1015 & ~n1016;
  assign n1018 = n155 & ~n1017;
  assign n1019 = ~n158 & ~n1018;
  assign n1020 = n157 & ~n1017;
  assign n1021 = n1019 & ~n1020;
  assign n1022 = n99 & ~n1021;
  assign n1023 = ~n100 & ~n1022;
  assign n1024 = n98 & ~n1021;
  assign n1025 = n1023 & ~n1024;
  assign n1026 = n96 & ~n1025;
  assign n1027 = n72 & n96;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = n72 & ~n1025;
  assign n1030 = n1028 & ~n1029;
  assign n1031 = n40 & ~n1030;
  assign n1032 = ~n43 & ~n1031;
  assign n1033 = n42 & ~n1030;
  assign n1034 = n1032 & ~n1033;
  assign n1035 = n23 & ~n1034;
  assign n1036 = ~n24 & ~n1035;
  assign n1037 = n22 & ~n1034;
  assign n1038 = n1036 & ~n1037;
  assign n1039 = n29 & ~n1038;
  assign n1040 = n25 & n29;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = n25 & ~n1038;
  assign n1043 = n1041 & ~n1042;
  assign n1044 = n304 & ~n361;
  assign n1045 = ~n364 & ~n1044;
  assign n1046 = n304 & ~n357;
  assign n1047 = n1045 & ~n1046;
  assign n1048 = ~n224 & n261;
  assign n1049 = n224 & ~n261;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = ~n263 & ~n1050;
  assign n1052 = n263 & n1050;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n1047 & ~n1053;
  assign n1055 = n226 & ~n1053;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = n226 & ~n1047;
  assign n1058 = n1056 & ~n1057;
  assign n1059 = ~n157 & ~n1017;
  assign n1060 = n157 & n1017;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = ~n155 & ~n1061;
  assign n1063 = n155 & n1061;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = ~n1058 & ~n1064;
  assign n1066 = n154 & ~n1064;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = n154 & ~n1058;
  assign n1069 = n1067 & ~n1068;
  assign n1070 = ~n98 & ~n1021;
  assign n1071 = n98 & n1021;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = ~n99 & ~n1072;
  assign n1074 = n99 & n1072;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = ~n1069 & ~n1075;
  assign n1077 = n126 & ~n1075;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n126 & ~n1069;
  assign n1080 = n1078 & ~n1079;
  assign n1081 = ~n72 & ~n1025;
  assign n1082 = n72 & n1025;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n96 & ~n1083;
  assign n1085 = n96 & n1083;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1080 & ~n1086;
  assign n1088 = n74 & ~n1086;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = n74 & ~n1080;
  assign n1091 = n1089 & ~n1090;
  assign n1092 = ~n42 & ~n1030;
  assign n1093 = n42 & n1030;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = ~n40 & ~n1094;
  assign n1096 = n40 & n1094;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = ~n1091 & ~n1097;
  assign n1099 = n39 & ~n1097;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = n39 & ~n1091;
  assign n1102 = n1100 & ~n1101;
  assign n1103 = ~n22 & ~n1034;
  assign n1104 = n22 & n1034;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = ~n23 & ~n1105;
  assign n1107 = n23 & n1105;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = ~n1102 & ~n1108;
  assign n1110 = n47 & ~n1108;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = n47 & ~n1102;
  assign n1113 = n1111 & ~n1112;
  assign n1114 = n400 & ~n460;
  assign n1115 = ~n463 & ~n1114;
  assign n1116 = n400 & ~n453;
  assign n1117 = n1115 & ~n1116;
  assign n1118 = ~n304 & ~n357;
  assign n1119 = n304 & n357;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = n361 & ~n1120;
  assign n1122 = ~n361 & n1120;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~n1117 & ~n1123;
  assign n1125 = n306 & ~n1123;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = n306 & ~n1117;
  assign n1128 = n1126 & ~n1127;
  assign n1129 = ~n226 & ~n1047;
  assign n1130 = n226 & n1047;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = n1053 & ~n1131;
  assign n1133 = ~n1053 & n1131;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n1128 & ~n1134;
  assign n1136 = n223 & ~n1134;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = n223 & ~n1128;
  assign n1139 = n1137 & ~n1138;
  assign n1140 = ~n154 & ~n1058;
  assign n1141 = n154 & n1058;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = n1064 & ~n1142;
  assign n1144 = ~n1064 & n1142;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = ~n1139 & ~n1145;
  assign n1147 = n192 & ~n1145;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = n192 & ~n1139;
  assign n1150 = n1148 & ~n1149;
  assign n1151 = ~n126 & ~n1069;
  assign n1152 = n126 & n1069;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = n1075 & ~n1153;
  assign n1155 = ~n1075 & n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = ~n1150 & ~n1156;
  assign n1158 = n128 & ~n1156;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = n128 & ~n1150;
  assign n1161 = n1159 & ~n1160;
  assign n1162 = ~n74 & ~n1080;
  assign n1163 = n74 & n1080;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = n1086 & ~n1164;
  assign n1166 = ~n1086 & n1164;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1161 & ~n1167;
  assign n1169 = n71 & ~n1167;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = n71 & ~n1161;
  assign n1172 = n1170 & ~n1171;
  assign n1173 = ~n39 & ~n1091;
  assign n1174 = n39 & n1091;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = n1097 & ~n1175;
  assign n1177 = ~n1097 & n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1172 & ~n1178;
  assign n1180 = n79 & ~n1178;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = n79 & ~n1172;
  assign n1183 = n1181 & ~n1182;
  assign n1184 = ~n400 & ~n453;
  assign n1185 = n400 & n453;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = n460 & ~n1186;
  assign n1188 = ~n460 & n1186;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = n499 & ~n551;
  assign n1191 = ~n560 & ~n1190;
  assign n1192 = n499 & ~n559;
  assign n1193 = n1191 & ~n1192;
  assign n1194 = ~n1189 & ~n1193;
  assign n1195 = n403 & ~n1189;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = n403 & ~n1193;
  assign n1198 = n1196 & ~n1197;
  assign n1199 = ~n306 & ~n1117;
  assign n1200 = n306 & n1117;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = n1123 & ~n1201;
  assign n1203 = ~n1123 & n1201;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~n1198 & ~n1204;
  assign n1206 = n303 & ~n1204;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = n303 & ~n1198;
  assign n1209 = n1207 & ~n1208;
  assign n1210 = ~n223 & ~n1128;
  assign n1211 = n223 & n1128;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = n1134 & ~n1212;
  assign n1214 = ~n1134 & n1212;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = ~n1209 & ~n1215;
  assign n1217 = n273 & ~n1215;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = n273 & ~n1209;
  assign n1220 = n1218 & ~n1219;
  assign n1221 = ~n192 & ~n1139;
  assign n1222 = n192 & n1139;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = n1145 & ~n1223;
  assign n1225 = ~n1145 & n1223;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = ~n1220 & ~n1226;
  assign n1228 = n194 & ~n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = n194 & ~n1220;
  assign n1231 = n1229 & ~n1230;
  assign n1232 = ~n128 & ~n1150;
  assign n1233 = n128 & n1150;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = n1156 & ~n1234;
  assign n1236 = ~n1156 & n1234;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~n1231 & ~n1237;
  assign n1239 = n125 & ~n1237;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = n125 & ~n1231;
  assign n1242 = n1240 & ~n1241;
  assign n1243 = ~n71 & ~n1161;
  assign n1244 = n71 & n1161;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = n1167 & ~n1245;
  assign n1247 = ~n1167 & n1245;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = ~n1242 & ~n1248;
  assign n1250 = n133 & ~n1248;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = n133 & ~n1242;
  assign n1253 = n1251 & ~n1252;
  assign n1254 = ~n403 & ~n1193;
  assign n1255 = n403 & n1193;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = n1189 & ~n1256;
  assign n1258 = ~n1189 & n1256;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n499 & ~n559;
  assign n1261 = n499 & n559;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = n551 & ~n1262;
  assign n1264 = ~n551 & n1262;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = n596 & ~n650;
  assign n1267 = ~n651 & ~n1266;
  assign n1268 = n596 & ~n644;
  assign n1269 = n1267 & ~n1268;
  assign n1270 = ~n1265 & ~n1269;
  assign n1271 = n502 & ~n1265;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = n502 & ~n1269;
  assign n1274 = n1272 & ~n1273;
  assign n1275 = ~n1259 & ~n1274;
  assign n1276 = n401 & ~n1259;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = n401 & ~n1274;
  assign n1279 = n1277 & ~n1278;
  assign n1280 = ~n303 & ~n1198;
  assign n1281 = n303 & n1198;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = n1204 & ~n1282;
  assign n1284 = ~n1204 & n1282;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~n1279 & ~n1285;
  assign n1287 = n370 & ~n1285;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = n370 & ~n1279;
  assign n1290 = n1288 & ~n1289;
  assign n1291 = ~n273 & ~n1209;
  assign n1292 = n273 & n1209;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n1215 & ~n1293;
  assign n1295 = ~n1215 & n1293;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~n1290 & ~n1296;
  assign n1298 = n275 & ~n1296;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = n275 & ~n1290;
  assign n1301 = n1299 & ~n1300;
  assign n1302 = ~n194 & ~n1220;
  assign n1303 = n194 & n1220;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n1226 & ~n1304;
  assign n1306 = ~n1226 & n1304;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1301 & ~n1307;
  assign n1309 = n191 & ~n1307;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = n191 & ~n1301;
  assign n1312 = n1310 & ~n1311;
  assign n1313 = ~n125 & ~n1231;
  assign n1314 = n125 & n1231;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = n1237 & ~n1315;
  assign n1317 = ~n1237 & n1315;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~n1312 & ~n1318;
  assign n1320 = n199 & ~n1318;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n199 & ~n1312;
  assign n1323 = n1321 & ~n1322;
  assign n1324 = ~n401 & ~n1274;
  assign n1325 = n401 & n1274;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = n1259 & ~n1326;
  assign n1328 = ~n1259 & n1326;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = ~n502 & ~n1269;
  assign n1331 = n502 & n1269;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = n1265 & ~n1332;
  assign n1334 = ~n1265 & n1332;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = n679 & ~n734;
  assign n1337 = ~n735 & ~n1336;
  assign n1338 = n679 & ~n728;
  assign n1339 = n1337 & ~n1338;
  assign n1340 = ~n596 & ~n644;
  assign n1341 = n596 & n644;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = n650 & ~n1342;
  assign n1344 = ~n650 & n1342;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1339 & ~n1345;
  assign n1347 = n598 & ~n1345;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = n598 & ~n1339;
  assign n1350 = n1348 & ~n1349;
  assign n1351 = ~n1335 & ~n1350;
  assign n1352 = n500 & ~n1335;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = n500 & ~n1350;
  assign n1355 = n1353 & ~n1354;
  assign n1356 = ~n1329 & ~n1355;
  assign n1357 = n468 & ~n1329;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = n468 & ~n1355;
  assign n1360 = n1358 & ~n1359;
  assign n1361 = ~n370 & ~n1279;
  assign n1362 = n370 & n1279;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1285 & ~n1363;
  assign n1365 = ~n1285 & n1363;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1360 & ~n1366;
  assign n1368 = n372 & ~n1366;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = n372 & ~n1360;
  assign n1371 = n1369 & ~n1370;
  assign n1372 = ~n275 & ~n1290;
  assign n1373 = n275 & n1290;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = n1296 & ~n1374;
  assign n1376 = ~n1296 & n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = ~n1371 & ~n1377;
  assign n1379 = n272 & ~n1377;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = n272 & ~n1371;
  assign n1382 = n1380 & ~n1381;
  assign n1383 = ~n191 & ~n1301;
  assign n1384 = n191 & n1301;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = n1307 & ~n1385;
  assign n1387 = ~n1307 & n1385;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = ~n1382 & ~n1388;
  assign n1390 = n268 & ~n1388;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = n268 & ~n1382;
  assign n1393 = n1391 & ~n1392;
  assign n1394 = ~n468 & ~n1355;
  assign n1395 = n468 & n1355;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = n1329 & ~n1396;
  assign n1398 = ~n1329 & n1396;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~n500 & ~n1350;
  assign n1401 = n500 & n1350;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = n1335 & ~n1402;
  assign n1404 = ~n1335 & n1402;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = n755 & ~n805;
  assign n1407 = ~n806 & ~n1406;
  assign n1408 = n755 & ~n799;
  assign n1409 = n1407 & ~n1408;
  assign n1410 = ~n679 & ~n728;
  assign n1411 = n679 & n728;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = n734 & ~n1412;
  assign n1414 = ~n734 & n1412;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~n1409 & ~n1415;
  assign n1417 = n681 & ~n1415;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = n681 & ~n1409;
  assign n1420 = n1418 & ~n1419;
  assign n1421 = ~n598 & ~n1339;
  assign n1422 = n598 & n1339;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = n1345 & ~n1423;
  assign n1425 = ~n1345 & n1423;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~n1420 & ~n1426;
  assign n1428 = n595 & ~n1426;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = n595 & ~n1420;
  assign n1431 = n1429 & ~n1430;
  assign n1432 = ~n1405 & ~n1431;
  assign n1433 = n565 & ~n1405;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = n565 & ~n1431;
  assign n1436 = n1434 & ~n1435;
  assign n1437 = ~n1399 & ~n1436;
  assign n1438 = n471 & ~n1399;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = n471 & ~n1436;
  assign n1441 = n1439 & ~n1440;
  assign n1442 = ~n372 & ~n1360;
  assign n1443 = n372 & n1360;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = n1366 & ~n1444;
  assign n1446 = ~n1366 & n1444;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1441 & ~n1447;
  assign n1449 = n369 & ~n1447;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = n369 & ~n1441;
  assign n1452 = n1450 & ~n1451;
  assign n1453 = ~n272 & ~n1371;
  assign n1454 = n272 & n1371;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = n1377 & ~n1455;
  assign n1457 = ~n1377 & n1455;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~n1452 & ~n1458;
  assign n1460 = n258 & ~n1458;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = n258 & ~n1452;
  assign n1463 = n1461 & ~n1462;
  assign n1464 = ~n471 & ~n1436;
  assign n1465 = n471 & n1436;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = n1399 & ~n1466;
  assign n1468 = ~n1399 & n1466;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = ~n565 & ~n1431;
  assign n1471 = n565 & n1431;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = n1405 & ~n1472;
  assign n1474 = ~n1405 & n1472;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n824 & ~n869;
  assign n1477 = ~n870 & ~n1476;
  assign n1478 = n824 & ~n863;
  assign n1479 = n1477 & ~n1478;
  assign n1480 = ~n755 & ~n799;
  assign n1481 = n755 & n799;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = n805 & ~n1482;
  assign n1484 = ~n805 & n1482;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~n1479 & ~n1485;
  assign n1487 = n757 & ~n1485;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = n757 & ~n1479;
  assign n1490 = n1488 & ~n1489;
  assign n1491 = ~n681 & ~n1409;
  assign n1492 = n681 & n1409;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = n1415 & ~n1493;
  assign n1495 = ~n1415 & n1493;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1490 & ~n1496;
  assign n1498 = n678 & ~n1496;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = n678 & ~n1490;
  assign n1501 = n1499 & ~n1500;
  assign n1502 = ~n595 & ~n1420;
  assign n1503 = n595 & n1420;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = n1426 & ~n1504;
  assign n1506 = ~n1426 & n1504;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1501 & ~n1507;
  assign n1509 = n656 & ~n1507;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = n656 & ~n1501;
  assign n1512 = n1510 & ~n1511;
  assign n1513 = ~n1475 & ~n1512;
  assign n1514 = n567 & ~n1475;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = n567 & ~n1512;
  assign n1517 = n1515 & ~n1516;
  assign n1518 = ~n1469 & ~n1517;
  assign n1519 = n469 & ~n1469;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = n469 & ~n1517;
  assign n1522 = n1520 & ~n1521;
  assign n1523 = ~n369 & ~n1441;
  assign n1524 = n369 & n1441;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = n1447 & ~n1525;
  assign n1527 = ~n1447 & n1525;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1522 & ~n1528;
  assign n1530 = n349 & ~n1528;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = n349 & ~n1522;
  assign n1533 = n1531 & ~n1532;
  assign n1534 = ~n913 & n955;
  assign n1535 = ~n914 & ~n1534;
  assign n1536 = ~n907 & n955;
  assign n1537 = n1535 & ~n1536;
  assign n1538 = ~n824 & ~n863;
  assign n1539 = n824 & n863;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = n869 & ~n1540;
  assign n1542 = ~n869 & n1540;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1537 & ~n1543;
  assign n1545 = n823 & ~n1543;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = n823 & ~n1537;
  assign n1548 = n1546 & ~n1547;
  assign n1549 = ~n757 & ~n1479;
  assign n1550 = n757 & n1479;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = n1485 & ~n1551;
  assign n1553 = ~n1485 & n1551;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~n1548 & ~n1554;
  assign n1556 = n754 & ~n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = n754 & ~n1548;
  assign n1559 = n1557 & ~n1558;
  assign n1560 = ~n678 & ~n1490;
  assign n1561 = n678 & n1490;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = n1496 & ~n1562;
  assign n1564 = ~n1496 & n1562;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~n1559 & ~n1565;
  assign n1567 = n752 & ~n1565;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = n752 & ~n1559;
  assign n1570 = n1568 & ~n1569;
  assign n1571 = ~n656 & ~n1501;
  assign n1572 = n656 & n1501;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = n1507 & ~n1573;
  assign n1575 = ~n1507 & n1573;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = ~n1570 & ~n1576;
  assign n1578 = n655 & ~n1576;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = n655 & ~n1570;
  assign n1581 = n1579 & ~n1580;
  assign n1582 = ~n567 & ~n1512;
  assign n1583 = n567 & n1512;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n1475 & ~n1584;
  assign n1586 = ~n1475 & n1584;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = ~n1581 & ~n1587;
  assign n1589 = n564 & ~n1587;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = n564 & ~n1581;
  assign n1592 = n1590 & ~n1591;
  assign n1593 = ~n469 & ~n1517;
  assign n1594 = n469 & n1517;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = n1469 & ~n1595;
  assign n1597 = ~n1469 & n1595;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1592 & ~n1598;
  assign n1600 = n445 & ~n1598;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = n445 & ~n1592;
  assign n1603 = n1601 & ~n1602;
  assign n1604 = ~n445 & ~n1592;
  assign n1605 = n445 & n1592;
  assign n1606 = ~n1604 & ~n1605;
  assign n1607 = n1598 & ~n1606;
  assign n1608 = ~n1598 & n1606;
  assign n1609 = ~n1607 & ~n1608;
  assign n1610 = ~n564 & ~n1581;
  assign n1611 = n564 & n1581;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = n1587 & ~n1612;
  assign n1614 = ~n1587 & n1612;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n655 & ~n1570;
  assign n1617 = n655 & n1570;
  assign n1618 = ~n1616 & ~n1617;
  assign n1619 = n1576 & ~n1618;
  assign n1620 = ~n1576 & n1618;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = ~n752 & ~n1559;
  assign n1623 = n752 & n1559;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = n1565 & ~n1624;
  assign n1626 = ~n1565 & n1624;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n754 & ~n1548;
  assign n1629 = n754 & n1548;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n1554 & ~n1630;
  assign n1632 = ~n1554 & n1630;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n823 & ~n1537;
  assign n1635 = n823 & n1537;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = n1543 & ~n1636;
  assign n1638 = ~n1543 & n1636;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = ~n907 & ~n955;
  assign n1641 = n907 & n955;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = n913 & ~n1642;
  assign n1644 = ~n913 & n1642;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = n951 & ~n1645;
  assign n1647 = ~n1639 & n1646;
  assign n1648 = ~n1633 & n1647;
  assign n1649 = ~n1627 & n1648;
  assign n1650 = ~n1621 & n1649;
  assign n1651 = ~n1615 & n1650;
  assign n1652 = ~n1609 & n1651;
  assign n1653 = ~n1603 & n1652;
  assign n1654 = ~n349 & ~n1522;
  assign n1655 = n349 & n1522;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = n1528 & ~n1656;
  assign n1658 = ~n1528 & n1656;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = n1652 & ~n1659;
  assign n1661 = ~n1653 & ~n1660;
  assign n1662 = ~n1603 & ~n1659;
  assign n1663 = n1661 & ~n1662;
  assign n1664 = ~n1533 & ~n1663;
  assign n1665 = ~n258 & ~n1452;
  assign n1666 = n258 & n1452;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = n1458 & ~n1667;
  assign n1669 = ~n1458 & n1667;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = ~n1663 & ~n1670;
  assign n1672 = ~n1664 & ~n1671;
  assign n1673 = ~n1533 & ~n1670;
  assign n1674 = n1672 & ~n1673;
  assign n1675 = ~n1463 & ~n1674;
  assign n1676 = ~n268 & ~n1382;
  assign n1677 = n268 & n1382;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = n1388 & ~n1678;
  assign n1680 = ~n1388 & n1678;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = ~n1674 & ~n1681;
  assign n1683 = ~n1675 & ~n1682;
  assign n1684 = ~n1463 & ~n1681;
  assign n1685 = n1683 & ~n1684;
  assign n1686 = ~n1393 & ~n1685;
  assign n1687 = ~n199 & ~n1312;
  assign n1688 = n199 & n1312;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = n1318 & ~n1689;
  assign n1691 = ~n1318 & n1689;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n1685 & ~n1692;
  assign n1694 = ~n1686 & ~n1693;
  assign n1695 = ~n1393 & ~n1692;
  assign n1696 = n1694 & ~n1695;
  assign n1697 = ~n1323 & ~n1696;
  assign n1698 = ~n133 & ~n1242;
  assign n1699 = n133 & n1242;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = n1248 & ~n1700;
  assign n1702 = ~n1248 & n1700;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = ~n1696 & ~n1703;
  assign n1705 = ~n1697 & ~n1704;
  assign n1706 = ~n1323 & ~n1703;
  assign n1707 = n1705 & ~n1706;
  assign n1708 = ~n1253 & ~n1707;
  assign n1709 = ~n79 & ~n1172;
  assign n1710 = n79 & n1172;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = n1178 & ~n1711;
  assign n1713 = ~n1178 & n1711;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~n1707 & ~n1714;
  assign n1716 = ~n1708 & ~n1715;
  assign n1717 = ~n1253 & ~n1714;
  assign n1718 = n1716 & ~n1717;
  assign n1719 = ~n1183 & ~n1718;
  assign n1720 = ~n47 & ~n1102;
  assign n1721 = n47 & n1102;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = n1108 & ~n1722;
  assign n1724 = ~n1108 & n1722;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = ~n1718 & ~n1725;
  assign n1727 = ~n1719 & ~n1726;
  assign n1728 = ~n1183 & ~n1725;
  assign n1729 = n1727 & ~n1728;
  assign n1730 = ~n1113 & ~n1729;
  assign n1731 = ~n25 & ~n1038;
  assign n1732 = n25 & n1038;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = ~n29 & ~n1733;
  assign n1735 = n29 & n1733;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = ~n1729 & ~n1736;
  assign n1738 = ~n1730 & ~n1737;
  assign n1739 = ~n1113 & ~n1736;
  assign n1740 = n1738 & ~n1739;
  assign n1741 = ~n1043 & ~n1740;
  assign n1742 = n31 & ~n1740;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = n31 & ~n1043;
  assign n1745 = n1743 & ~n1744;
  assign n1746 = ~n1013 & n1745;
  assign n1747 = n1013 & ~n1745;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = n183 & ~n996;
  assign n1750 = n1001 & ~n1749;
  assign n1751 = n38 & ~n63;
  assign n1752 = ~n38 & n63;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1750 & n1753;
  assign n1755 = n1750 & ~n1753;
  assign n1756 = ~n1754 & ~n1755;
  assign n1757 = ~n31 & ~n1043;
  assign n1758 = n31 & n1043;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = n1740 & ~n1759;
  assign n1761 = ~n1740 & n1759;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~n1756 & n1762;
  assign n1764 = n1756 & ~n1762;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~n182 & ~n996;
  assign n1767 = ~n998 & ~n1766;
  assign n1768 = n70 & ~n117;
  assign n1769 = ~n70 & n117;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~n1767 & n1770;
  assign n1772 = n1767 & ~n1770;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = ~n1113 & n1736;
  assign n1775 = n1113 & ~n1736;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n1729 & ~n1776;
  assign n1778 = ~n1729 & n1776;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = ~n1773 & n1779;
  assign n1781 = n1773 & ~n1779;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = n124 & ~n181;
  assign n1784 = ~n124 & n181;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = ~n996 & n1785;
  assign n1787 = n996 & ~n1785;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = ~n1183 & n1725;
  assign n1790 = n1183 & ~n1725;
  assign n1791 = ~n1789 & ~n1790;
  assign n1792 = n1718 & ~n1791;
  assign n1793 = ~n1718 & n1791;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = ~n1788 & n1794;
  assign n1796 = n1788 & ~n1794;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~n335 & n532;
  assign n1799 = n845 & n1798;
  assign n1800 = ~n972 & n1799;
  assign n1801 = ~n983 & n1798;
  assign n1802 = ~n335 & ~n988;
  assign n1803 = ~n990 & ~n1802;
  assign n1804 = ~n1801 & n1803;
  assign n1805 = ~n1800 & n1804;
  assign n1806 = n190 & ~n250;
  assign n1807 = ~n190 & n250;
  assign n1808 = ~n1806 & ~n1807;
  assign n1809 = ~n1805 & n1808;
  assign n1810 = n1805 & ~n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~n1253 & n1714;
  assign n1813 = n1253 & ~n1714;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = n1707 & ~n1814;
  assign n1816 = ~n1707 & n1814;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = ~n1811 & n1817;
  assign n1819 = n1811 & ~n1817;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = n532 & n845;
  assign n1822 = ~n972 & n1821;
  assign n1823 = n532 & ~n983;
  assign n1824 = n988 & ~n1823;
  assign n1825 = ~n1822 & n1824;
  assign n1826 = n257 & ~n334;
  assign n1827 = ~n257 & n334;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1825 & n1828;
  assign n1830 = n1825 & ~n1828;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1323 & n1703;
  assign n1833 = n1323 & ~n1703;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = n1696 & ~n1834;
  assign n1836 = ~n1696 & n1834;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1831 & n1837;
  assign n1839 = n1831 & ~n1837;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n531 & n845;
  assign n1842 = ~n972 & n1841;
  assign n1843 = ~n531 & ~n983;
  assign n1844 = ~n985 & ~n1843;
  assign n1845 = ~n1842 & n1844;
  assign n1846 = n342 & ~n431;
  assign n1847 = ~n342 & n431;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~n1845 & n1848;
  assign n1850 = n1845 & ~n1848;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = ~n1393 & n1692;
  assign n1853 = n1393 & ~n1692;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = n1685 & ~n1854;
  assign n1856 = ~n1685 & n1854;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~n1851 & n1857;
  assign n1859 = n1851 & ~n1857;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = n845 & ~n972;
  assign n1862 = n983 & ~n1861;
  assign n1863 = n438 & ~n530;
  assign n1864 = ~n438 & n530;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1862 & n1865;
  assign n1867 = n1862 & ~n1865;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = ~n1463 & n1681;
  assign n1870 = n1463 & ~n1681;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = n1674 & ~n1871;
  assign n1873 = ~n1674 & n1871;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1868 & n1874;
  assign n1876 = n1868 & ~n1874;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = ~n710 & n844;
  assign n1879 = ~n972 & n1878;
  assign n1880 = ~n710 & ~n977;
  assign n1881 = ~n979 & ~n1880;
  assign n1882 = ~n1879 & n1881;
  assign n1883 = n539 & ~n626;
  assign n1884 = ~n539 & n626;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = ~n1882 & n1885;
  assign n1887 = n1882 & ~n1885;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = ~n1533 & n1670;
  assign n1890 = n1533 & ~n1670;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = n1663 & ~n1891;
  assign n1893 = ~n1663 & n1891;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = ~n1888 & n1894;
  assign n1896 = n1888 & ~n1894;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = n844 & ~n972;
  assign n1899 = n977 & ~n1898;
  assign n1900 = n633 & ~n709;
  assign n1901 = ~n633 & n709;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = ~n1899 & n1902;
  assign n1904 = n1899 & ~n1902;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1603 & n1659;
  assign n1907 = n1603 & ~n1659;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~n1652 & ~n1908;
  assign n1910 = n1652 & n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n1905 & n1911;
  assign n1913 = n1905 & ~n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n843 & ~n972;
  assign n1916 = ~n974 & ~n1915;
  assign n1917 = n717 & ~n781;
  assign n1918 = ~n717 & n781;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = ~n1916 & n1919;
  assign n1921 = n1916 & ~n1919;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = n1609 & n1651;
  assign n1924 = ~n1609 & ~n1651;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = ~n1922 & n1925;
  assign n1927 = n1922 & ~n1925;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = n788 & ~n842;
  assign n1930 = ~n788 & n842;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = ~n972 & n1931;
  assign n1933 = n972 & ~n1931;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1615 & n1650;
  assign n1936 = ~n1615 & ~n1650;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = ~n1934 & n1937;
  assign n1939 = n1934 & ~n1937;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~n931 & n966;
  assign n1942 = ~n968 & ~n1941;
  assign n1943 = n852 & ~n889;
  assign n1944 = ~n852 & n889;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = ~n1942 & n1945;
  assign n1947 = n1942 & ~n1945;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = n1621 & n1649;
  assign n1950 = ~n1621 & ~n1649;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = ~n1948 & n1951;
  assign n1953 = n1948 & ~n1951;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = n896 & ~n930;
  assign n1956 = ~n896 & n930;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = n966 & n1957;
  assign n1959 = ~n966 & ~n1957;
  assign n1960 = ~n1958 & ~n1959;
  assign n1961 = n1627 & n1648;
  assign n1962 = ~n1627 & ~n1648;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = ~n1960 & n1963;
  assign n1965 = n1960 & ~n1963;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = n938 & ~n965;
  assign n1968 = ~n938 & n965;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = n1633 & n1647;
  assign n1971 = ~n1633 & ~n1647;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1969 & n1972;
  assign n1974 = n1969 & ~n1972;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = n956 & n961;
  assign n1977 = ~n956 & ~n961;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n957 & ~n1978;
  assign n1980 = n957 & n1978;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = n1639 & n1646;
  assign n1983 = ~n1639 & ~n1646;
  assign n1984 = ~n1982 & ~n1983;
  assign n1985 = ~n1981 & n1984;
  assign n1986 = n1981 & ~n1984;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = ~n954 & ~n955;
  assign n1989 = n954 & n955;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = n951 & n1645;
  assign n1992 = ~n951 & ~n1645;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n1990 & n1993;
  assign n1995 = n1990 & ~n1993;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = n1987 & n1996;
  assign n1998 = n1975 & n1997;
  assign n1999 = n1966 & n1998;
  assign n2000 = n1954 & n1999;
  assign n2001 = n1940 & n2000;
  assign n2002 = n1928 & n2001;
  assign n2003 = n1914 & n2002;
  assign n2004 = n1897 & n2003;
  assign n2005 = n1877 & n2004;
  assign n2006 = n1860 & n2005;
  assign n2007 = n1840 & n2006;
  assign n2008 = n1820 & n2007;
  assign n2009 = n1797 & n2008;
  assign n2010 = n1782 & n2009;
  assign n2011 = n1765 & n2010;
  assign po0 = ~n1748 | ~n2011;
endmodule


