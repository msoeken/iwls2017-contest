// Benchmark "" written by ABC on Wed Apr 26 17:08:30 2017

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107;
  wire n316, n317, n319, n320, n321, n322, n323, n324, n326, n327, n328,
    n329, n330, n331, n333, n334, n335, n336, n337, n338, n340, n341, n342,
    n343, n344, n345, n348, n349, n350, n351, n352, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1958,
    n1959, n1960, n1961, n1962, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2002,
    n2003, n2004, n2005, n2006, n2008, n2009, n2010, n2011, n2012, n2013,
    n2015, n2016, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
    n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2520, n2521, n2523, n2524, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2558, n2559, n2560, n2561, n2562, n2564,
    n2565, n2566, n2567, n2568, n2569, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2591, n2592, n2593, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2607, n2608,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2639, n2640, n2642,
    n2643, n2644, n2645, n2646, n2647, n2649, n2650, n2651, n2652, n2653,
    n2655, n2656, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2671, n2672, n2673, n2674, n2675, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2699, n2700, n2701, n2702, n2703, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2716, n2717, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2730, n2731, n2733,
    n2734, n2735, n2736, n2737, n2738, n2740, n2741, n2742, n2743, n2744,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207;
  assign n316 = ~pi001 & ~pi020;
  assign n317 = pi001 & pi020;
  assign po041 = ~n316 | n317;
  assign n319 = pi107 & pi163;
  assign n320 = pi073 & ~pi107;
  assign n321 = pi073 & pi151;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~pi107 & pi151;
  assign n324 = n322 & ~n323;
  assign po042 = ~n319 | n324;
  assign n326 = pi133 & pi153;
  assign n327 = pi075 & ~pi133;
  assign n328 = pi075 & pi141;
  assign n329 = ~n327 & ~n328;
  assign n330 = ~pi133 & pi141;
  assign n331 = n329 & ~n330;
  assign po043 = ~n326 | n331;
  assign n333 = pi106 & pi109;
  assign n334 = pi105 & ~pi106;
  assign n335 = pi105 & pi108;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~pi106 & pi108;
  assign n338 = n336 & ~n337;
  assign po044 = ~n333 | n338;
  assign n340 = pi095 & pi122;
  assign n341 = pi085 & ~pi095;
  assign n342 = pi085 & pi111;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~pi095 & pi111;
  assign n345 = n343 & ~n344;
  assign po045 = ~n340 | n345;
  assign po048 = pi001 | ~pi165;
  assign n348 = pi001 & pi066;
  assign n349 = pi001 & ~pi067;
  assign n350 = ~n348 & ~n349;
  assign n351 = pi066 & ~pi067;
  assign n352 = n350 & ~n351;
  assign po051 = ~pi066 | ~n352;
  assign po055 = pi000 & pi086;
  assign n355 = pi005 & pi012;
  assign n356 = pi005 & pi186;
  assign n357 = ~n355 & ~n356;
  assign n358 = pi012 & pi186;
  assign n359 = n357 & ~n358;
  assign n360 = pi012 & n359;
  assign n361 = ~pi005 & ~pi012;
  assign n362 = ~n355 & n361;
  assign n363 = pi186 & n362;
  assign n364 = ~n360 & ~n363;
  assign n365 = n360 & n363;
  assign n366 = n364 & ~n365;
  assign n367 = ~pi205 & ~n366;
  assign n368 = pi205 & n366;
  assign po056 = ~n367 & ~n368;
  assign n370 = pi173 & ~pi206;
  assign n371 = pi011 & n370;
  assign n372 = pi172 & pi173;
  assign n373 = pi172 & n370;
  assign n374 = ~n372 & ~n373;
  assign n375 = pi173 & n370;
  assign n376 = n374 & ~n375;
  assign n377 = pi011 & n376;
  assign n378 = ~n371 & ~n377;
  assign n379 = n370 & n376;
  assign n380 = n378 & ~n379;
  assign n381 = pi002 & pi003;
  assign n382 = pi005 & n381;
  assign n383 = pi005 & ~pi136;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~pi136 & n381;
  assign n386 = n384 & ~n385;
  assign n387 = ~n381 & n386;
  assign n388 = n381 & ~n386;
  assign n389 = n387 & ~n388;
  assign n390 = ~pi171 & ~n389;
  assign n391 = pi171 & n389;
  assign n392 = ~n390 & ~n391;
  assign n393 = pi005 & ~pi137;
  assign n394 = ~n382 & ~n393;
  assign n395 = ~pi137 & n381;
  assign n396 = n394 & ~n395;
  assign n397 = ~n381 & n396;
  assign n398 = n381 & ~n396;
  assign n399 = n397 & ~n398;
  assign n400 = ~pi170 & ~n399;
  assign n401 = pi170 & n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n392 & n402;
  assign n404 = pi005 & ~pi138;
  assign n405 = ~n382 & ~n404;
  assign n406 = ~pi138 & n381;
  assign n407 = n405 & ~n406;
  assign n408 = ~n381 & n407;
  assign n409 = n381 & ~n407;
  assign n410 = n408 & ~n409;
  assign n411 = pi053 & ~n410;
  assign n412 = ~pi168 & ~n381;
  assign n413 = pi168 & n381;
  assign n414 = n412 & ~n413;
  assign n415 = pi005 & ~pi132;
  assign n416 = ~n382 & ~n415;
  assign n417 = ~pi132 & n381;
  assign n418 = n416 & ~n417;
  assign n419 = n414 & n418;
  assign n420 = ~n414 & ~n418;
  assign n421 = n419 & ~n420;
  assign n422 = pi005 & ~pi139;
  assign n423 = ~n382 & ~n422;
  assign n424 = ~pi139 & n381;
  assign n425 = n423 & ~n424;
  assign n426 = ~n381 & n425;
  assign n427 = n381 & ~n425;
  assign n428 = n426 & ~n427;
  assign n429 = ~pi169 & ~n428;
  assign n430 = pi169 & n428;
  assign n431 = ~n429 & ~n430;
  assign n432 = n421 & ~n431;
  assign n433 = pi053 & ~n432;
  assign n434 = ~n411 & ~n433;
  assign n435 = ~n410 & ~n432;
  assign n436 = n434 & ~n435;
  assign n437 = ~n392 & ~n436;
  assign n438 = ~n403 & ~n437;
  assign n439 = n402 & ~n436;
  assign n440 = n438 & ~n439;
  assign n441 = ~n392 & n440;
  assign n442 = pi171 & ~n389;
  assign n443 = ~pi170 & n399;
  assign n444 = pi170 & ~n399;
  assign n445 = n443 & ~n444;
  assign n446 = pi171 & ~n445;
  assign n447 = ~n442 & ~n446;
  assign n448 = ~n389 & ~n445;
  assign n449 = n447 & ~n448;
  assign n450 = ~n441 & ~n449;
  assign n451 = ~pi053 & ~n410;
  assign n452 = pi053 & n410;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~pi005 & ~pi132;
  assign n455 = pi005 & pi132;
  assign n456 = n454 & ~n455;
  assign n457 = ~pi132 & ~n456;
  assign n458 = ~n417 & ~n457;
  assign n459 = n381 & ~n456;
  assign n460 = n458 & ~n459;
  assign n461 = ~pi168 & ~n460;
  assign n462 = pi168 & n460;
  assign n463 = ~n461 & ~n462;
  assign n464 = n453 & ~n463;
  assign n465 = ~n431 & ~n463;
  assign n466 = ~n464 & ~n465;
  assign n467 = ~n431 & n453;
  assign n468 = n466 & ~n467;
  assign n469 = ~n453 & ~n468;
  assign n470 = ~n402 & n469;
  assign n471 = pi005 & ~pi077;
  assign n472 = ~n382 & ~n471;
  assign n473 = ~pi077 & n381;
  assign n474 = n472 & ~n473;
  assign n475 = ~n381 & n474;
  assign n476 = n381 & ~n474;
  assign n477 = n475 & ~n476;
  assign n478 = ~pi183 & ~n477;
  assign n479 = pi183 & n477;
  assign n480 = ~n478 & ~n479;
  assign n481 = pi005 & ~pi078;
  assign n482 = ~n382 & ~n481;
  assign n483 = ~pi078 & n381;
  assign n484 = n482 & ~n483;
  assign n485 = ~n381 & n484;
  assign n486 = n381 & ~n484;
  assign n487 = n485 & ~n486;
  assign n488 = ~pi182 & ~n487;
  assign n489 = pi182 & n487;
  assign n490 = ~n488 & ~n489;
  assign n491 = pi005 & ~pi079;
  assign n492 = ~n382 & ~n491;
  assign n493 = ~pi079 & n381;
  assign n494 = n492 & ~n493;
  assign n495 = ~n381 & n494;
  assign n496 = n381 & ~n494;
  assign n497 = n495 & ~n496;
  assign n498 = ~pi181 & ~n497;
  assign n499 = pi181 & n497;
  assign n500 = ~n498 & ~n499;
  assign n501 = ~n490 & ~n500;
  assign n502 = n480 & n501;
  assign n503 = pi005 & ~pi076;
  assign n504 = ~n382 & ~n503;
  assign n505 = ~pi076 & n381;
  assign n506 = n504 & ~n505;
  assign n507 = ~n381 & n506;
  assign n508 = n381 & ~n506;
  assign n509 = n507 & ~n508;
  assign n510 = ~pi184 & ~n509;
  assign n511 = pi184 & n509;
  assign n512 = ~n510 & ~n511;
  assign n513 = n480 & ~n512;
  assign n514 = ~n502 & ~n513;
  assign n515 = n501 & ~n512;
  assign n516 = n514 & ~n515;
  assign n517 = ~n480 & ~n516;
  assign n518 = pi005 & ~pi080;
  assign n519 = ~n382 & ~n518;
  assign n520 = ~pi080 & n381;
  assign n521 = n519 & ~n520;
  assign n522 = ~n381 & n521;
  assign n523 = n381 & ~n521;
  assign n524 = n522 & ~n523;
  assign n525 = pi180 & ~n524;
  assign n526 = pi068 & pi081;
  assign n527 = ~pi005 & pi081;
  assign n528 = pi005 & ~pi081;
  assign n529 = ~n527 & ~n528;
  assign n530 = pi068 & n529;
  assign n531 = ~n526 & ~n530;
  assign n532 = pi081 & n529;
  assign n533 = n531 & ~n532;
  assign n534 = ~pi179 & ~n533;
  assign n535 = pi071 & pi082;
  assign n536 = ~pi005 & pi082;
  assign n537 = pi005 & ~pi082;
  assign n538 = ~n536 & ~n537;
  assign n539 = pi071 & n538;
  assign n540 = ~n535 & ~n539;
  assign n541 = pi082 & n538;
  assign n542 = n540 & ~n541;
  assign n543 = ~pi178 & ~n542;
  assign n544 = pi069 & pi083;
  assign n545 = ~pi005 & pi083;
  assign n546 = pi005 & ~pi083;
  assign n547 = ~n545 & ~n546;
  assign n548 = pi069 & n547;
  assign n549 = ~n544 & ~n548;
  assign n550 = pi083 & n547;
  assign n551 = n549 & ~n550;
  assign n552 = ~pi177 & ~n551;
  assign n553 = pi177 & n551;
  assign n554 = ~n552 & ~n553;
  assign n555 = pi072 & pi074;
  assign n556 = ~pi005 & pi074;
  assign n557 = pi005 & ~pi074;
  assign n558 = ~n556 & ~n557;
  assign n559 = pi072 & n558;
  assign n560 = ~n555 & ~n559;
  assign n561 = pi074 & n558;
  assign n562 = n560 & ~n561;
  assign n563 = ~pi176 & ~n562;
  assign n564 = n554 & n563;
  assign n565 = ~n552 & ~n564;
  assign n566 = n552 & n564;
  assign n567 = n565 & ~n566;
  assign n568 = ~pi178 & ~n567;
  assign n569 = ~n543 & ~n568;
  assign n570 = ~n542 & ~n567;
  assign n571 = n569 & ~n570;
  assign n572 = ~pi179 & ~n571;
  assign n573 = ~n534 & ~n572;
  assign n574 = ~n533 & ~n571;
  assign n575 = n573 & ~n574;
  assign n576 = pi180 & n575;
  assign n577 = ~n525 & ~n576;
  assign n578 = ~n524 & n575;
  assign n579 = n577 & ~n578;
  assign n580 = n517 & n579;
  assign n581 = pi184 & ~n509;
  assign n582 = pi183 & ~n477;
  assign n583 = pi182 & ~n487;
  assign n584 = ~pi181 & n497;
  assign n585 = pi181 & ~n497;
  assign n586 = n584 & ~n585;
  assign n587 = pi182 & ~n586;
  assign n588 = ~n583 & ~n587;
  assign n589 = ~n487 & ~n586;
  assign n590 = n588 & ~n589;
  assign n591 = pi183 & ~n590;
  assign n592 = ~n582 & ~n591;
  assign n593 = ~n477 & ~n590;
  assign n594 = n592 & ~n593;
  assign n595 = pi184 & ~n594;
  assign n596 = ~n581 & ~n595;
  assign n597 = ~n509 & ~n594;
  assign n598 = n596 & ~n597;
  assign n599 = ~n580 & ~n598;
  assign n600 = pi009 & pi144;
  assign n601 = ~pi005 & pi144;
  assign n602 = pi005 & ~pi144;
  assign n603 = ~n601 & ~n602;
  assign n604 = pi009 & n603;
  assign n605 = ~n600 & ~n604;
  assign n606 = pi144 & n603;
  assign n607 = n605 & ~n606;
  assign n608 = ~pi202 & ~n607;
  assign n609 = pi202 & n607;
  assign n610 = ~n608 & ~n609;
  assign n611 = pi010 & pi145;
  assign n612 = ~pi005 & pi145;
  assign n613 = pi005 & ~pi145;
  assign n614 = ~n612 & ~n613;
  assign n615 = pi010 & n614;
  assign n616 = ~n611 & ~n615;
  assign n617 = pi145 & n614;
  assign n618 = n616 & ~n617;
  assign n619 = ~pi201 & ~n618;
  assign n620 = pi201 & n618;
  assign n621 = ~n619 & ~n620;
  assign n622 = n610 & n621;
  assign n623 = ~n610 & ~n621;
  assign n624 = n622 & ~n623;
  assign n625 = pi015 & pi143;
  assign n626 = ~pi005 & pi143;
  assign n627 = pi005 & ~pi143;
  assign n628 = ~n626 & ~n627;
  assign n629 = pi015 & n628;
  assign n630 = ~n625 & ~n629;
  assign n631 = pi143 & n628;
  assign n632 = n630 & ~n631;
  assign n633 = ~pi203 & ~n632;
  assign n634 = pi203 & n632;
  assign n635 = ~n633 & ~n634;
  assign n636 = n624 & n635;
  assign n637 = ~n624 & ~n635;
  assign n638 = n636 & ~n637;
  assign n639 = pi014 & pi146;
  assign n640 = ~pi005 & pi146;
  assign n641 = pi005 & ~pi146;
  assign n642 = ~n640 & ~n641;
  assign n643 = pi014 & n642;
  assign n644 = ~n639 & ~n643;
  assign n645 = pi146 & n642;
  assign n646 = n644 & ~n645;
  assign n647 = ~pi200 & ~n646;
  assign n648 = pi200 & n646;
  assign n649 = ~n647 & ~n648;
  assign n650 = pi062 & pi147;
  assign n651 = ~pi005 & pi147;
  assign n652 = pi005 & ~pi147;
  assign n653 = ~n651 & ~n652;
  assign n654 = pi062 & n653;
  assign n655 = ~n650 & ~n654;
  assign n656 = pi147 & n653;
  assign n657 = n655 & ~n656;
  assign n658 = ~pi199 & ~n657;
  assign n659 = pi199 & n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n649 & n660;
  assign n662 = pi049 & pi148;
  assign n663 = ~pi005 & pi148;
  assign n664 = pi005 & ~pi148;
  assign n665 = ~n663 & ~n664;
  assign n666 = pi049 & n665;
  assign n667 = ~n662 & ~n666;
  assign n668 = pi148 & n665;
  assign n669 = n667 & ~n668;
  assign n670 = ~pi198 & ~n669;
  assign n671 = pi061 & pi140;
  assign n672 = ~pi005 & pi140;
  assign n673 = pi005 & ~pi140;
  assign n674 = ~n672 & ~n673;
  assign n675 = pi061 & n674;
  assign n676 = ~n671 & ~n675;
  assign n677 = pi140 & n674;
  assign n678 = n676 & ~n677;
  assign n679 = ~pi196 & ~n678;
  assign n680 = pi050 & pi149;
  assign n681 = ~pi005 & pi149;
  assign n682 = pi005 & ~pi149;
  assign n683 = ~n681 & ~n682;
  assign n684 = pi050 & n683;
  assign n685 = ~n680 & ~n684;
  assign n686 = pi149 & n683;
  assign n687 = n685 & ~n686;
  assign n688 = ~pi197 & ~n687;
  assign n689 = pi197 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = n679 & n690;
  assign n692 = ~pi198 & n691;
  assign n693 = ~n670 & ~n692;
  assign n694 = ~n669 & n691;
  assign n695 = n693 & ~n694;
  assign n696 = ~n649 & ~n695;
  assign n697 = ~n661 & ~n696;
  assign n698 = n660 & ~n695;
  assign n699 = n697 & ~n698;
  assign n700 = n649 & ~n699;
  assign n701 = ~pi200 & n658;
  assign n702 = ~n647 & ~n701;
  assign n703 = ~n646 & n658;
  assign n704 = n702 & ~n703;
  assign n705 = ~n700 & n704;
  assign n706 = n700 & ~n704;
  assign n707 = n705 & ~n706;
  assign n708 = pi198 & n669;
  assign n709 = ~n670 & ~n708;
  assign n710 = pi196 & n678;
  assign n711 = ~n679 & ~n710;
  assign n712 = n709 & ~n711;
  assign n713 = ~n690 & ~n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n690 & n709;
  assign n716 = n714 & ~n715;
  assign n717 = n709 & n716;
  assign n718 = ~n709 & ~n716;
  assign n719 = n717 & ~n718;
  assign n720 = n660 & n719;
  assign n721 = ~n660 & ~n719;
  assign n722 = n720 & ~n721;
  assign n723 = pi051 & pi154;
  assign n724 = ~pi005 & pi154;
  assign n725 = pi005 & ~pi154;
  assign n726 = ~n724 & ~n725;
  assign n727 = pi051 & n726;
  assign n728 = ~n723 & ~n727;
  assign n729 = pi154 & n726;
  assign n730 = n728 & ~n729;
  assign n731 = ~pi194 & ~n730;
  assign n732 = pi194 & n730;
  assign n733 = ~n731 & ~n732;
  assign n734 = pi063 & pi155;
  assign n735 = ~pi005 & pi155;
  assign n736 = pi005 & ~pi155;
  assign n737 = ~n735 & ~n736;
  assign n738 = pi063 & n737;
  assign n739 = ~n734 & ~n738;
  assign n740 = pi155 & n737;
  assign n741 = n739 & ~n740;
  assign n742 = ~pi193 & ~n741;
  assign n743 = pi193 & n741;
  assign n744 = ~n742 & ~n743;
  assign n745 = n733 & n744;
  assign n746 = ~n733 & ~n744;
  assign n747 = n745 & ~n746;
  assign n748 = pi064 & pi156;
  assign n749 = ~pi005 & pi156;
  assign n750 = pi005 & ~pi156;
  assign n751 = ~n749 & ~n750;
  assign n752 = pi064 & n751;
  assign n753 = ~n748 & ~n752;
  assign n754 = pi156 & n751;
  assign n755 = n753 & ~n754;
  assign n756 = ~pi192 & ~n755;
  assign n757 = pi065 & pi157;
  assign n758 = ~pi005 & pi157;
  assign n759 = pi005 & ~pi157;
  assign n760 = ~n758 & ~n759;
  assign n761 = pi065 & n760;
  assign n762 = ~n757 & ~n761;
  assign n763 = pi157 & n760;
  assign n764 = n762 & ~n763;
  assign n765 = ~pi191 & ~n764;
  assign n766 = ~pi192 & n765;
  assign n767 = ~n756 & ~n766;
  assign n768 = ~n755 & n765;
  assign n769 = n767 & ~n768;
  assign n770 = n747 & ~n769;
  assign n771 = ~pi194 & n742;
  assign n772 = ~n731 & ~n771;
  assign n773 = ~n730 & n742;
  assign n774 = n772 & ~n773;
  assign n775 = ~n770 & n774;
  assign n776 = n770 & ~n774;
  assign n777 = n775 & ~n776;
  assign n778 = pi052 & pi158;
  assign n779 = ~pi005 & pi158;
  assign n780 = pi005 & ~pi158;
  assign n781 = ~n779 & ~n780;
  assign n782 = pi052 & n781;
  assign n783 = ~n778 & ~n782;
  assign n784 = pi158 & n781;
  assign n785 = n783 & ~n784;
  assign n786 = pi190 & n785;
  assign n787 = pi006 & pi159;
  assign n788 = ~pi005 & pi159;
  assign n789 = pi005 & ~pi159;
  assign n790 = ~n788 & ~n789;
  assign n791 = pi006 & n790;
  assign n792 = ~n787 & ~n791;
  assign n793 = pi159 & n790;
  assign n794 = n792 & ~n793;
  assign n795 = pi189 & n794;
  assign n796 = ~pi189 & ~n794;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n786 & n797;
  assign n799 = n786 & ~n797;
  assign n800 = n798 & ~n799;
  assign n801 = pi007 & pi160;
  assign n802 = ~pi005 & pi160;
  assign n803 = pi005 & ~pi160;
  assign n804 = ~n802 & ~n803;
  assign n805 = pi007 & n804;
  assign n806 = ~n801 & ~n805;
  assign n807 = pi160 & n804;
  assign n808 = n806 & ~n807;
  assign n809 = ~pi188 & ~n808;
  assign n810 = pi188 & n808;
  assign n811 = ~n809 & ~n810;
  assign n812 = n786 & n811;
  assign n813 = pi008 & pi161;
  assign n814 = ~pi005 & pi161;
  assign n815 = pi005 & ~pi161;
  assign n816 = ~n814 & ~n815;
  assign n817 = pi008 & n816;
  assign n818 = ~n813 & ~n817;
  assign n819 = pi161 & n816;
  assign n820 = n818 & ~n819;
  assign n821 = ~pi187 & ~n820;
  assign n822 = pi187 & n820;
  assign n823 = ~n821 & ~n822;
  assign n824 = pi205 & ~n823;
  assign n825 = ~n368 & ~n824;
  assign n826 = n366 & ~n823;
  assign n827 = n825 & ~n826;
  assign n828 = n823 & ~n827;
  assign n829 = n786 & n828;
  assign n830 = ~n812 & ~n829;
  assign n831 = n811 & n828;
  assign n832 = n830 & ~n831;
  assign n833 = n800 & ~n832;
  assign n834 = ~pi190 & ~n785;
  assign n835 = n360 & n823;
  assign n836 = ~n821 & ~n835;
  assign n837 = n821 & n835;
  assign n838 = n836 & ~n837;
  assign n839 = ~pi188 & ~n838;
  assign n840 = ~n809 & ~n839;
  assign n841 = ~n808 & ~n838;
  assign n842 = n840 & ~n841;
  assign n843 = ~pi189 & ~n842;
  assign n844 = ~n796 & ~n843;
  assign n845 = ~n794 & ~n842;
  assign n846 = n844 & ~n845;
  assign n847 = ~pi190 & ~n846;
  assign n848 = ~n834 & ~n847;
  assign n849 = ~n785 & ~n846;
  assign n850 = n848 & ~n849;
  assign n851 = ~n833 & n850;
  assign n852 = n833 & ~n850;
  assign n853 = n851 & ~n852;
  assign n854 = pi192 & n755;
  assign n855 = ~n756 & ~n854;
  assign n856 = pi191 & n764;
  assign n857 = ~n765 & ~n856;
  assign n858 = n855 & ~n857;
  assign n859 = ~n747 & n855;
  assign n860 = ~n858 & ~n859;
  assign n861 = ~n747 & ~n857;
  assign n862 = n860 & ~n861;
  assign n863 = n855 & n862;
  assign n864 = ~n855 & ~n862;
  assign n865 = n863 & ~n864;
  assign n866 = ~n853 & n865;
  assign n867 = ~n774 & ~n853;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n774 & n865;
  assign n870 = n868 & ~n869;
  assign n871 = n777 & n870;
  assign n872 = ~n777 & ~n870;
  assign n873 = n871 & ~n872;
  assign n874 = n649 & ~n873;
  assign n875 = ~n719 & ~n873;
  assign n876 = ~n874 & ~n875;
  assign n877 = n649 & ~n719;
  assign n878 = n876 & ~n877;
  assign n879 = n722 & ~n878;
  assign n880 = ~n700 & n879;
  assign n881 = n660 & n688;
  assign n882 = ~n649 & ~n709;
  assign n883 = ~n661 & ~n882;
  assign n884 = n660 & ~n709;
  assign n885 = n883 & ~n884;
  assign n886 = n881 & n885;
  assign n887 = n879 & n886;
  assign n888 = ~n880 & ~n887;
  assign n889 = ~n700 & n886;
  assign n890 = n888 & ~n889;
  assign n891 = n707 & n890;
  assign n892 = ~n707 & ~n890;
  assign n893 = n891 & ~n892;
  assign n894 = ~n624 & ~n893;
  assign n895 = pi029 & pi142;
  assign n896 = ~pi005 & pi142;
  assign n897 = pi005 & ~pi142;
  assign n898 = ~n896 & ~n897;
  assign n899 = pi029 & n898;
  assign n900 = ~n895 & ~n899;
  assign n901 = pi142 & n898;
  assign n902 = n900 & ~n901;
  assign n903 = ~pi204 & ~n902;
  assign n904 = pi204 & n902;
  assign n905 = ~n903 & ~n904;
  assign n906 = ~n893 & n905;
  assign n907 = ~n894 & ~n906;
  assign n908 = ~n624 & n905;
  assign n909 = n907 & ~n908;
  assign n910 = n638 & ~n909;
  assign n911 = ~pi202 & n619;
  assign n912 = ~n608 & ~n911;
  assign n913 = ~n607 & n619;
  assign n914 = n912 & ~n913;
  assign n915 = ~pi203 & ~n914;
  assign n916 = ~n633 & ~n915;
  assign n917 = ~n632 & ~n914;
  assign n918 = n916 & ~n917;
  assign n919 = ~pi204 & ~n918;
  assign n920 = ~n903 & ~n919;
  assign n921 = ~n902 & ~n918;
  assign n922 = n920 & ~n921;
  assign n923 = ~n910 & n922;
  assign n924 = n910 & ~n922;
  assign n925 = n923 & ~n924;
  assign n926 = ~pi180 & ~n524;
  assign n927 = pi180 & n524;
  assign n928 = ~n926 & ~n927;
  assign n929 = pi179 & n533;
  assign n930 = ~n534 & ~n929;
  assign n931 = pi178 & n542;
  assign n932 = ~n543 & ~n931;
  assign n933 = n554 & ~n932;
  assign n934 = pi176 & n562;
  assign n935 = ~n563 & ~n934;
  assign n936 = ~n932 & ~n935;
  assign n937 = ~n933 & ~n936;
  assign n938 = n554 & ~n935;
  assign n939 = n937 & ~n938;
  assign n940 = n554 & n939;
  assign n941 = ~n554 & ~n939;
  assign n942 = n940 & ~n941;
  assign n943 = n930 & n942;
  assign n944 = ~n930 & ~n942;
  assign n945 = n943 & ~n944;
  assign n946 = ~n928 & n945;
  assign n947 = n517 & n946;
  assign n948 = ~n925 & n947;
  assign n949 = n580 & ~n925;
  assign n950 = ~n948 & ~n949;
  assign n951 = n580 & n947;
  assign n952 = n950 & ~n951;
  assign n953 = n599 & n952;
  assign n954 = n392 & n953;
  assign n955 = n469 & n953;
  assign n956 = ~n954 & ~n955;
  assign n957 = n392 & n469;
  assign n958 = n956 & ~n957;
  assign n959 = n470 & n958;
  assign n960 = ~n441 & n959;
  assign n961 = ~pi169 & n428;
  assign n962 = pi169 & ~n428;
  assign n963 = n961 & ~n962;
  assign n964 = ~n402 & n963;
  assign n965 = ~n392 & ~n453;
  assign n966 = ~n403 & ~n965;
  assign n967 = n402 & ~n453;
  assign n968 = n966 & ~n967;
  assign n969 = n964 & ~n968;
  assign n970 = n959 & n969;
  assign n971 = ~n960 & ~n970;
  assign n972 = ~n441 & n969;
  assign n973 = n971 & ~n972;
  assign n974 = n450 & n973;
  assign n975 = n380 & n974;
  assign n976 = ~pi011 & pi172;
  assign n977 = ~pi011 & pi173;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n372 & n978;
  assign n980 = pi206 & ~n979;
  assign n981 = ~pi011 & n980;
  assign n982 = pi011 & ~n980;
  assign n983 = ~n981 & ~n982;
  assign n984 = n380 & ~n983;
  assign n985 = ~n975 & ~n984;
  assign n986 = n974 & ~n983;
  assign n987 = n985 & ~n986;
  assign po057 = ~n380 | n987;
  assign n989 = ~pi011 & pi206;
  assign n990 = pi166 & pi174;
  assign n991 = pi011 & pi166;
  assign n992 = pi011 & pi174;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n990 & n993;
  assign n995 = n989 & n994;
  assign n996 = pi005 & ~pi090;
  assign n997 = ~n382 & ~n996;
  assign n998 = ~pi090 & n381;
  assign n999 = n997 & ~n998;
  assign n1000 = ~n381 & n999;
  assign n1001 = n381 & ~n999;
  assign n1002 = n1000 & ~n1001;
  assign n1003 = pi057 & ~pi170;
  assign n1004 = ~pi005 & pi057;
  assign n1005 = pi005 & ~pi057;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = pi057 & ~n1006;
  assign n1008 = ~n1003 & ~n1007;
  assign n1009 = ~pi170 & ~n1006;
  assign n1010 = n1008 & ~n1009;
  assign n1011 = ~n1002 & n1010;
  assign n1012 = pi056 & ~pi169;
  assign n1013 = ~pi005 & pi056;
  assign n1014 = pi005 & ~pi056;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = pi056 & ~n1015;
  assign n1017 = ~n1012 & ~n1016;
  assign n1018 = ~pi169 & ~n1015;
  assign n1019 = n1017 & ~n1018;
  assign n1020 = pi005 & pi092;
  assign n1021 = pi005 & ~n1020;
  assign n1022 = ~n382 & ~n1021;
  assign n1023 = n381 & ~n1020;
  assign n1024 = n1022 & ~n1023;
  assign n1025 = n1019 & ~n1024;
  assign n1026 = ~n1019 & n1024;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = ~n1011 & n1027;
  assign n1029 = n1011 & ~n1027;
  assign n1030 = n1028 & ~n1029;
  assign n1031 = n1002 & n1010;
  assign n1032 = ~n1002 & ~n1010;
  assign n1033 = n1031 & ~n1032;
  assign n1034 = n1002 & ~n1033;
  assign n1035 = pi005 & ~pi091;
  assign n1036 = ~n382 & ~n1035;
  assign n1037 = ~pi091 & n381;
  assign n1038 = n1036 & ~n1037;
  assign n1039 = ~n381 & n1038;
  assign n1040 = n381 & ~n1038;
  assign n1041 = n1039 & ~n1040;
  assign n1042 = pi046 & ~pi053;
  assign n1043 = ~pi005 & pi046;
  assign n1044 = pi005 & ~pi046;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = pi046 & ~n1045;
  assign n1047 = ~n1042 & ~n1046;
  assign n1048 = ~pi053 & ~n1045;
  assign n1049 = n1047 & ~n1048;
  assign n1050 = n1041 & ~n1049;
  assign n1051 = n1002 & n1050;
  assign n1052 = ~n1034 & ~n1051;
  assign n1053 = ~n1033 & n1050;
  assign n1054 = n1052 & ~n1053;
  assign n1055 = ~n1011 & ~n1054;
  assign n1056 = ~n1041 & n1049;
  assign n1057 = ~n1054 & n1056;
  assign n1058 = ~n1055 & ~n1057;
  assign n1059 = ~n1011 & n1056;
  assign n1060 = n1058 & ~n1059;
  assign n1061 = n1030 & n1060;
  assign n1062 = ~n1030 & ~n1060;
  assign n1063 = n1061 & ~n1062;
  assign n1064 = pi005 & ~pi096;
  assign n1065 = ~n382 & ~n1064;
  assign n1066 = ~pi096 & n381;
  assign n1067 = n1065 & ~n1066;
  assign n1068 = ~n381 & n1067;
  assign n1069 = n381 & ~n1067;
  assign n1070 = n1068 & ~n1069;
  assign n1071 = pi055 & ~pi184;
  assign n1072 = ~pi005 & pi055;
  assign n1073 = pi005 & ~pi055;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = pi055 & ~n1074;
  assign n1076 = ~n1071 & ~n1075;
  assign n1077 = ~pi184 & ~n1074;
  assign n1078 = n1076 & ~n1077;
  assign n1079 = n1070 & ~n1078;
  assign n1080 = ~n1070 & n1078;
  assign n1081 = pi005 & ~pi097;
  assign n1082 = ~n382 & ~n1081;
  assign n1083 = ~pi097 & n381;
  assign n1084 = n1082 & ~n1083;
  assign n1085 = ~n381 & n1084;
  assign n1086 = n381 & ~n1084;
  assign n1087 = n1085 & ~n1086;
  assign n1088 = pi054 & ~pi183;
  assign n1089 = ~pi005 & pi054;
  assign n1090 = pi005 & ~pi054;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = pi054 & ~n1091;
  assign n1093 = ~n1088 & ~n1092;
  assign n1094 = ~pi183 & ~n1091;
  assign n1095 = n1093 & ~n1094;
  assign n1096 = n1087 & ~n1095;
  assign n1097 = pi005 & ~pi098;
  assign n1098 = ~n382 & ~n1097;
  assign n1099 = ~pi098 & n381;
  assign n1100 = n1098 & ~n1099;
  assign n1101 = ~n381 & n1100;
  assign n1102 = n381 & ~n1100;
  assign n1103 = n1101 & ~n1102;
  assign n1104 = pi045 & ~pi182;
  assign n1105 = ~pi005 & pi045;
  assign n1106 = pi005 & ~pi045;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = pi045 & ~n1107;
  assign n1109 = ~n1104 & ~n1108;
  assign n1110 = ~pi182 & ~n1107;
  assign n1111 = n1109 & ~n1110;
  assign n1112 = n1103 & ~n1111;
  assign n1113 = n1087 & n1112;
  assign n1114 = ~n1096 & ~n1113;
  assign n1115 = ~n1095 & n1112;
  assign n1116 = n1114 & ~n1115;
  assign n1117 = ~n1080 & ~n1116;
  assign n1118 = ~n1079 & ~n1117;
  assign n1119 = n1079 & n1117;
  assign n1120 = n1118 & ~n1119;
  assign n1121 = ~n1103 & n1111;
  assign n1122 = ~n1112 & ~n1121;
  assign n1123 = ~n1087 & n1095;
  assign n1124 = ~n1096 & ~n1123;
  assign n1125 = n1122 & n1124;
  assign n1126 = ~n1122 & ~n1124;
  assign n1127 = n1125 & ~n1126;
  assign n1128 = pi005 & ~pi099;
  assign n1129 = ~n382 & ~n1128;
  assign n1130 = ~pi099 & n381;
  assign n1131 = n1129 & ~n1130;
  assign n1132 = ~n381 & n1131;
  assign n1133 = n381 & ~n1131;
  assign n1134 = n1132 & ~n1133;
  assign n1135 = pi026 & ~pi181;
  assign n1136 = ~pi005 & pi026;
  assign n1137 = pi005 & ~pi026;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = pi026 & ~n1138;
  assign n1140 = ~n1135 & ~n1139;
  assign n1141 = ~pi181 & ~n1138;
  assign n1142 = n1140 & ~n1141;
  assign n1143 = ~n1134 & ~n1142;
  assign n1144 = ~n1079 & ~n1080;
  assign n1145 = ~n1134 & n1144;
  assign n1146 = ~n1143 & ~n1145;
  assign n1147 = ~n1142 & n1144;
  assign n1148 = n1146 & ~n1147;
  assign n1149 = n1134 & ~n1148;
  assign n1150 = ~pi005 & pi180;
  assign n1151 = pi005 & ~pi100;
  assign n1152 = ~n382 & ~n1151;
  assign n1153 = ~pi100 & n381;
  assign n1154 = n1152 & ~n1153;
  assign n1155 = ~n381 & n1154;
  assign n1156 = n381 & ~n1154;
  assign n1157 = n1155 & ~n1156;
  assign n1158 = ~pi005 & ~n1157;
  assign n1159 = ~n1150 & ~n1158;
  assign n1160 = pi180 & ~n1157;
  assign n1161 = n1159 & ~n1160;
  assign n1162 = pi005 & ~pi027;
  assign n1163 = pi005 & ~n1157;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = ~pi027 & ~n1157;
  assign n1166 = n1164 & ~n1165;
  assign n1167 = ~n1161 & ~n1166;
  assign n1168 = pi005 & pi180;
  assign n1169 = ~n1163 & ~n1168;
  assign n1170 = ~n1160 & n1169;
  assign n1171 = pi005 & pi027;
  assign n1172 = pi005 & n1157;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = pi027 & n1157;
  assign n1175 = n1173 & ~n1174;
  assign n1176 = n1170 & ~n1175;
  assign n1177 = pi068 & pi101;
  assign n1178 = ~pi005 & pi101;
  assign n1179 = pi005 & ~pi101;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = pi068 & n1180;
  assign n1182 = ~n1177 & ~n1181;
  assign n1183 = pi101 & n1180;
  assign n1184 = n1182 & ~n1183;
  assign n1185 = pi044 & ~pi179;
  assign n1186 = ~pi005 & pi044;
  assign n1187 = pi005 & ~pi044;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = pi044 & ~n1188;
  assign n1190 = ~n1185 & ~n1189;
  assign n1191 = ~pi179 & ~n1188;
  assign n1192 = n1190 & ~n1191;
  assign n1193 = n1184 & n1192;
  assign n1194 = ~n1184 & ~n1192;
  assign n1195 = n1193 & ~n1194;
  assign n1196 = pi071 & pi102;
  assign n1197 = ~pi005 & pi102;
  assign n1198 = pi005 & ~pi102;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = pi071 & n1199;
  assign n1201 = ~n1196 & ~n1200;
  assign n1202 = pi102 & n1199;
  assign n1203 = n1201 & ~n1202;
  assign n1204 = pi043 & ~pi178;
  assign n1205 = ~pi005 & pi043;
  assign n1206 = pi005 & ~pi043;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = pi043 & ~n1207;
  assign n1209 = ~n1204 & ~n1208;
  assign n1210 = ~pi178 & ~n1207;
  assign n1211 = n1209 & ~n1210;
  assign n1212 = ~n1203 & ~n1211;
  assign n1213 = pi069 & pi103;
  assign n1214 = ~pi005 & pi103;
  assign n1215 = pi005 & ~pi103;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = pi069 & n1216;
  assign n1218 = ~n1213 & ~n1217;
  assign n1219 = pi103 & n1216;
  assign n1220 = n1218 & ~n1219;
  assign n1221 = pi042 & ~pi177;
  assign n1222 = ~pi005 & pi042;
  assign n1223 = pi005 & ~pi042;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = pi042 & ~n1224;
  assign n1226 = ~n1221 & ~n1225;
  assign n1227 = ~pi177 & ~n1224;
  assign n1228 = n1226 & ~n1227;
  assign n1229 = ~n1220 & ~n1228;
  assign n1230 = pi072 & pi094;
  assign n1231 = ~pi005 & pi094;
  assign n1232 = pi005 & ~pi094;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = pi072 & n1233;
  assign n1235 = ~n1230 & ~n1234;
  assign n1236 = pi094 & n1233;
  assign n1237 = n1235 & ~n1236;
  assign n1238 = pi028 & ~pi176;
  assign n1239 = ~pi005 & pi028;
  assign n1240 = pi005 & ~pi028;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = pi028 & ~n1241;
  assign n1243 = ~n1238 & ~n1242;
  assign n1244 = ~pi176 & ~n1241;
  assign n1245 = n1243 & ~n1244;
  assign n1246 = ~n1237 & ~n1245;
  assign n1247 = ~n1220 & n1246;
  assign n1248 = ~n1229 & ~n1247;
  assign n1249 = ~n1228 & n1246;
  assign n1250 = n1248 & ~n1249;
  assign n1251 = ~n1212 & n1250;
  assign n1252 = n1212 & ~n1250;
  assign n1253 = n1251 & ~n1252;
  assign n1254 = ~n1195 & ~n1253;
  assign n1255 = ~n1195 & ~n1203;
  assign n1256 = ~n1212 & ~n1255;
  assign n1257 = ~n1195 & ~n1211;
  assign n1258 = n1256 & ~n1257;
  assign n1259 = n1254 & ~n1258;
  assign n1260 = ~n1176 & ~n1259;
  assign n1261 = n1176 & n1259;
  assign n1262 = n1260 & ~n1261;
  assign n1263 = n1176 & ~n1184;
  assign n1264 = ~n1194 & ~n1263;
  assign n1265 = n1176 & ~n1192;
  assign n1266 = n1264 & ~n1265;
  assign n1267 = n1262 & n1266;
  assign n1268 = ~n1262 & ~n1266;
  assign n1269 = n1267 & ~n1268;
  assign n1270 = n1167 & ~n1269;
  assign n1271 = n1149 & ~n1270;
  assign n1272 = n1134 & ~n1142;
  assign n1273 = ~n1134 & n1142;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = n1144 & n1274;
  assign n1276 = ~n1144 & ~n1274;
  assign n1277 = n1275 & ~n1276;
  assign n1278 = ~n1269 & n1277;
  assign n1279 = n1270 & n1277;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~n1269 & n1270;
  assign n1282 = n1280 & ~n1281;
  assign n1283 = n1149 & ~n1282;
  assign n1284 = ~n1271 & ~n1283;
  assign n1285 = ~n1270 & ~n1282;
  assign n1286 = n1284 & ~n1285;
  assign n1287 = n1127 & ~n1286;
  assign n1288 = n1117 & n1127;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = n1117 & ~n1286;
  assign n1291 = n1289 & ~n1290;
  assign n1292 = n1120 & n1291;
  assign n1293 = ~n1120 & ~n1291;
  assign n1294 = n1292 & ~n1293;
  assign n1295 = pi029 & pi112;
  assign n1296 = ~pi005 & pi112;
  assign n1297 = pi005 & ~pi112;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = pi029 & n1298;
  assign n1300 = ~n1295 & ~n1299;
  assign n1301 = pi112 & n1298;
  assign n1302 = n1300 & ~n1301;
  assign n1303 = pi025 & ~pi204;
  assign n1304 = ~pi005 & pi025;
  assign n1305 = pi005 & ~pi025;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = pi025 & ~n1306;
  assign n1308 = ~n1303 & ~n1307;
  assign n1309 = ~pi204 & ~n1306;
  assign n1310 = n1308 & ~n1309;
  assign n1311 = n1302 & n1310;
  assign n1312 = ~n1302 & ~n1310;
  assign n1313 = n1311 & ~n1312;
  assign n1314 = pi015 & pi113;
  assign n1315 = ~pi005 & pi113;
  assign n1316 = pi005 & ~pi113;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = pi015 & n1317;
  assign n1319 = ~n1314 & ~n1318;
  assign n1320 = pi113 & n1317;
  assign n1321 = n1319 & ~n1320;
  assign n1322 = pi024 & ~pi203;
  assign n1323 = ~pi005 & pi024;
  assign n1324 = pi005 & ~pi024;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = pi024 & ~n1325;
  assign n1327 = ~n1322 & ~n1326;
  assign n1328 = ~pi203 & ~n1325;
  assign n1329 = n1327 & ~n1328;
  assign n1330 = ~n1321 & ~n1329;
  assign n1331 = pi009 & pi114;
  assign n1332 = ~pi005 & pi114;
  assign n1333 = pi005 & ~pi114;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = pi009 & n1334;
  assign n1336 = ~n1331 & ~n1335;
  assign n1337 = pi114 & n1334;
  assign n1338 = n1336 & ~n1337;
  assign n1339 = pi023 & ~pi202;
  assign n1340 = ~pi005 & pi023;
  assign n1341 = pi005 & ~pi023;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = pi023 & ~n1342;
  assign n1344 = ~n1339 & ~n1343;
  assign n1345 = ~pi202 & ~n1342;
  assign n1346 = n1344 & ~n1345;
  assign n1347 = ~n1338 & ~n1346;
  assign n1348 = ~n1321 & n1347;
  assign n1349 = ~n1330 & ~n1348;
  assign n1350 = ~n1329 & n1347;
  assign n1351 = n1349 & ~n1350;
  assign n1352 = ~n1313 & ~n1351;
  assign n1353 = pi038 & ~pi201;
  assign n1354 = ~pi005 & pi038;
  assign n1355 = pi005 & ~pi038;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = pi038 & ~n1356;
  assign n1358 = ~n1353 & ~n1357;
  assign n1359 = ~pi201 & ~n1356;
  assign n1360 = n1358 & ~n1359;
  assign n1361 = n1338 & ~n1346;
  assign n1362 = ~n1338 & n1346;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1321 & ~n1329;
  assign n1365 = ~n1321 & n1329;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1363 & ~n1366;
  assign n1368 = ~n1360 & n1367;
  assign n1369 = n1302 & ~n1310;
  assign n1370 = ~n1302 & n1310;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~n1367 & ~n1371;
  assign n1373 = pi010 & pi115;
  assign n1374 = ~pi005 & pi115;
  assign n1375 = pi005 & ~pi115;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = pi010 & n1376;
  assign n1378 = ~n1373 & ~n1377;
  assign n1379 = pi115 & n1376;
  assign n1380 = n1378 & ~n1379;
  assign n1381 = ~n1371 & ~n1380;
  assign n1382 = ~n1372 & ~n1381;
  assign n1383 = ~n1367 & ~n1380;
  assign n1384 = n1382 & ~n1383;
  assign n1385 = n1368 & ~n1384;
  assign n1386 = ~n1352 & ~n1385;
  assign n1387 = n1352 & n1385;
  assign n1388 = n1386 & ~n1387;
  assign n1389 = ~n1302 & n1385;
  assign n1390 = ~n1312 & ~n1389;
  assign n1391 = ~n1310 & n1385;
  assign n1392 = n1390 & ~n1391;
  assign n1393 = n1388 & n1392;
  assign n1394 = ~n1388 & ~n1392;
  assign n1395 = n1393 & ~n1394;
  assign n1396 = ~n1360 & n1380;
  assign n1397 = n1360 & ~n1380;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n1371 & ~n1398;
  assign n1400 = ~n1372 & ~n1399;
  assign n1401 = ~n1367 & ~n1398;
  assign n1402 = n1400 & ~n1401;
  assign n1403 = n1367 & ~n1402;
  assign n1404 = pi014 & pi116;
  assign n1405 = ~pi005 & pi116;
  assign n1406 = pi005 & ~pi116;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = pi014 & n1407;
  assign n1409 = ~n1404 & ~n1408;
  assign n1410 = pi116 & n1407;
  assign n1411 = n1409 & ~n1410;
  assign n1412 = pi039 & ~pi200;
  assign n1413 = ~pi005 & pi039;
  assign n1414 = pi005 & ~pi039;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = pi039 & ~n1415;
  assign n1417 = ~n1412 & ~n1416;
  assign n1418 = ~pi200 & ~n1415;
  assign n1419 = n1417 & ~n1418;
  assign n1420 = ~n1411 & ~n1419;
  assign n1421 = pi062 & pi117;
  assign n1422 = ~pi005 & pi117;
  assign n1423 = pi005 & ~pi117;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = pi062 & n1424;
  assign n1426 = ~n1421 & ~n1425;
  assign n1427 = pi117 & n1424;
  assign n1428 = n1426 & ~n1427;
  assign n1429 = pi040 & ~pi199;
  assign n1430 = ~pi005 & pi040;
  assign n1431 = pi005 & ~pi040;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = pi040 & ~n1432;
  assign n1434 = ~n1429 & ~n1433;
  assign n1435 = ~pi199 & ~n1432;
  assign n1436 = n1434 & ~n1435;
  assign n1437 = ~n1428 & ~n1436;
  assign n1438 = pi049 & pi118;
  assign n1439 = ~pi005 & pi118;
  assign n1440 = pi005 & ~pi118;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = pi049 & n1441;
  assign n1443 = ~n1438 & ~n1442;
  assign n1444 = pi118 & n1441;
  assign n1445 = n1443 & ~n1444;
  assign n1446 = pi022 & ~pi198;
  assign n1447 = ~pi005 & pi022;
  assign n1448 = pi005 & ~pi022;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = pi022 & ~n1449;
  assign n1451 = ~n1446 & ~n1450;
  assign n1452 = ~pi198 & ~n1449;
  assign n1453 = n1451 & ~n1452;
  assign n1454 = ~n1445 & ~n1453;
  assign n1455 = pi005 & pi050;
  assign n1456 = pi037 & ~pi197;
  assign n1457 = ~pi005 & pi037;
  assign n1458 = pi005 & ~pi037;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = pi037 & ~n1459;
  assign n1461 = ~n1456 & ~n1460;
  assign n1462 = ~pi197 & ~n1459;
  assign n1463 = n1461 & ~n1462;
  assign n1464 = pi005 & ~n1463;
  assign n1465 = ~n1455 & ~n1464;
  assign n1466 = pi050 & ~n1463;
  assign n1467 = n1465 & ~n1466;
  assign n1468 = ~pi005 & pi119;
  assign n1469 = ~pi005 & ~n1463;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = pi119 & ~n1463;
  assign n1472 = n1470 & ~n1471;
  assign n1473 = ~n1467 & ~n1472;
  assign n1474 = pi061 & pi110;
  assign n1475 = ~pi005 & pi110;
  assign n1476 = pi005 & ~pi110;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = pi061 & n1477;
  assign n1479 = ~n1474 & ~n1478;
  assign n1480 = pi110 & n1477;
  assign n1481 = n1479 & ~n1480;
  assign n1482 = pi036 & ~pi196;
  assign n1483 = ~pi005 & pi036;
  assign n1484 = pi005 & ~pi036;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = pi036 & ~n1485;
  assign n1487 = ~n1482 & ~n1486;
  assign n1488 = ~pi196 & ~n1485;
  assign n1489 = n1487 & ~n1488;
  assign n1490 = ~n1481 & ~n1489;
  assign n1491 = n1473 & ~n1481;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = n1473 & ~n1489;
  assign n1494 = n1492 & ~n1493;
  assign n1495 = ~n1473 & n1494;
  assign n1496 = n1473 & ~n1494;
  assign n1497 = n1495 & ~n1496;
  assign n1498 = ~pi005 & pi050;
  assign n1499 = ~n1469 & ~n1498;
  assign n1500 = ~n1466 & n1499;
  assign n1501 = pi005 & pi119;
  assign n1502 = ~n1464 & ~n1501;
  assign n1503 = ~n1471 & n1502;
  assign n1504 = n1500 & n1503;
  assign n1505 = ~n1500 & ~n1503;
  assign n1506 = n1504 & ~n1505;
  assign n1507 = ~n1497 & ~n1506;
  assign n1508 = ~n1445 & n1507;
  assign n1509 = ~n1454 & ~n1508;
  assign n1510 = ~n1453 & n1507;
  assign n1511 = n1509 & ~n1510;
  assign n1512 = ~n1437 & n1511;
  assign n1513 = n1437 & ~n1511;
  assign n1514 = n1512 & ~n1513;
  assign n1515 = n1420 & ~n1514;
  assign n1516 = ~n1428 & n1436;
  assign n1517 = ~n1436 & n1516;
  assign n1518 = n1411 & n1419;
  assign n1519 = ~n1420 & n1518;
  assign n1520 = ~n1436 & ~n1519;
  assign n1521 = ~n1517 & ~n1520;
  assign n1522 = n1516 & ~n1519;
  assign n1523 = n1521 & ~n1522;
  assign n1524 = ~n1514 & n1523;
  assign n1525 = n1420 & ~n1524;
  assign n1526 = ~n1515 & ~n1525;
  assign n1527 = ~n1514 & ~n1524;
  assign n1528 = n1526 & ~n1527;
  assign n1529 = n1403 & ~n1528;
  assign n1530 = ~n1395 & n1403;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~n1395 & ~n1528;
  assign n1533 = n1531 & ~n1532;
  assign n1534 = n1395 & n1533;
  assign n1535 = ~n1395 & ~n1533;
  assign n1536 = n1534 & ~n1535;
  assign n1537 = pi063 & pi124;
  assign n1538 = ~pi005 & pi124;
  assign n1539 = pi005 & ~pi124;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = pi063 & n1540;
  assign n1542 = ~n1537 & ~n1541;
  assign n1543 = pi124 & n1540;
  assign n1544 = n1542 & ~n1543;
  assign n1545 = pi018 & ~pi193;
  assign n1546 = ~pi005 & pi018;
  assign n1547 = pi005 & ~pi018;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = pi018 & ~n1548;
  assign n1550 = ~n1545 & ~n1549;
  assign n1551 = ~pi193 & ~n1548;
  assign n1552 = n1550 & ~n1551;
  assign n1553 = n1544 & ~n1552;
  assign n1554 = ~n1544 & n1552;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = pi051 & pi123;
  assign n1557 = ~pi005 & pi123;
  assign n1558 = pi005 & ~pi123;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = pi051 & n1559;
  assign n1561 = ~n1556 & ~n1560;
  assign n1562 = pi123 & n1559;
  assign n1563 = n1561 & ~n1562;
  assign n1564 = pi019 & ~pi194;
  assign n1565 = ~pi005 & pi019;
  assign n1566 = pi005 & ~pi019;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = pi019 & ~n1567;
  assign n1569 = ~n1564 & ~n1568;
  assign n1570 = ~pi194 & ~n1567;
  assign n1571 = n1569 & ~n1570;
  assign n1572 = n1563 & ~n1571;
  assign n1573 = ~n1563 & n1571;
  assign n1574 = ~n1572 & ~n1573;
  assign n1575 = ~n1555 & ~n1574;
  assign n1576 = pi064 & pi125;
  assign n1577 = ~pi005 & pi125;
  assign n1578 = pi005 & ~pi125;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = pi064 & n1579;
  assign n1581 = ~n1576 & ~n1580;
  assign n1582 = pi125 & n1579;
  assign n1583 = n1581 & ~n1582;
  assign n1584 = pi017 & ~pi192;
  assign n1585 = ~pi005 & pi017;
  assign n1586 = pi005 & ~pi017;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = pi017 & ~n1587;
  assign n1589 = ~n1584 & ~n1588;
  assign n1590 = ~pi192 & ~n1587;
  assign n1591 = n1589 & ~n1590;
  assign n1592 = ~n1583 & ~n1591;
  assign n1593 = pi065 & pi126;
  assign n1594 = ~pi005 & pi126;
  assign n1595 = pi005 & ~pi126;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = pi065 & n1596;
  assign n1598 = ~n1593 & ~n1597;
  assign n1599 = pi126 & n1596;
  assign n1600 = n1598 & ~n1599;
  assign n1601 = pi016 & ~pi191;
  assign n1602 = ~pi005 & pi016;
  assign n1603 = pi005 & ~pi016;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = pi016 & ~n1604;
  assign n1606 = ~n1601 & ~n1605;
  assign n1607 = ~pi191 & ~n1604;
  assign n1608 = n1606 & ~n1607;
  assign n1609 = ~n1600 & ~n1608;
  assign n1610 = ~n1583 & n1609;
  assign n1611 = ~n1592 & ~n1610;
  assign n1612 = ~n1591 & n1609;
  assign n1613 = n1611 & ~n1612;
  assign n1614 = n1575 & ~n1613;
  assign n1615 = ~n1563 & ~n1571;
  assign n1616 = ~n1544 & ~n1552;
  assign n1617 = ~n1563 & n1616;
  assign n1618 = ~n1615 & ~n1617;
  assign n1619 = ~n1571 & n1616;
  assign n1620 = n1618 & ~n1619;
  assign n1621 = ~n1614 & ~n1620;
  assign n1622 = n1600 & ~n1608;
  assign n1623 = ~n1600 & n1608;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = n1583 & ~n1591;
  assign n1626 = ~n1583 & n1591;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n1624 & ~n1627;
  assign n1629 = n1575 & n1628;
  assign n1630 = pi052 & pi127;
  assign n1631 = ~pi005 & pi127;
  assign n1632 = pi005 & ~pi127;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = pi052 & n1633;
  assign n1635 = ~n1630 & ~n1634;
  assign n1636 = pi127 & n1633;
  assign n1637 = n1635 & ~n1636;
  assign n1638 = pi032 & ~pi190;
  assign n1639 = ~pi005 & pi032;
  assign n1640 = pi005 & ~pi032;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = pi032 & ~n1641;
  assign n1643 = ~n1638 & ~n1642;
  assign n1644 = ~pi190 & ~n1641;
  assign n1645 = n1643 & ~n1644;
  assign n1646 = n1637 & n1645;
  assign n1647 = ~n1637 & ~n1645;
  assign n1648 = n1646 & ~n1647;
  assign n1649 = pi006 & pi128;
  assign n1650 = ~pi005 & pi128;
  assign n1651 = pi005 & ~pi128;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = pi006 & n1652;
  assign n1654 = ~n1649 & ~n1653;
  assign n1655 = pi128 & n1652;
  assign n1656 = n1654 & ~n1655;
  assign n1657 = pi034 & ~pi189;
  assign n1658 = ~pi005 & pi034;
  assign n1659 = pi005 & ~pi034;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = pi034 & ~n1660;
  assign n1662 = ~n1657 & ~n1661;
  assign n1663 = ~pi189 & ~n1660;
  assign n1664 = n1662 & ~n1663;
  assign n1665 = ~n1656 & ~n1664;
  assign n1666 = pi007 & pi129;
  assign n1667 = ~pi005 & pi129;
  assign n1668 = pi005 & ~pi129;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = pi007 & n1669;
  assign n1671 = ~n1666 & ~n1670;
  assign n1672 = pi129 & n1669;
  assign n1673 = n1671 & ~n1672;
  assign n1674 = pi035 & ~pi188;
  assign n1675 = ~pi005 & pi035;
  assign n1676 = pi005 & ~pi035;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = pi035 & ~n1677;
  assign n1679 = ~n1674 & ~n1678;
  assign n1680 = ~pi188 & ~n1677;
  assign n1681 = n1679 & ~n1680;
  assign n1682 = n1673 & n1681;
  assign n1683 = ~n1673 & ~n1681;
  assign n1684 = n1682 & ~n1683;
  assign n1685 = ~pi005 & pi031;
  assign n1686 = pi033 & ~pi187;
  assign n1687 = ~pi005 & pi033;
  assign n1688 = pi005 & ~pi033;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = pi033 & ~n1689;
  assign n1691 = ~n1686 & ~n1690;
  assign n1692 = ~pi187 & ~n1689;
  assign n1693 = n1691 & ~n1692;
  assign n1694 = pi008 & ~n1693;
  assign n1695 = ~pi005 & ~n1693;
  assign n1696 = ~pi005 & pi008;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = ~n1694 & n1697;
  assign n1699 = pi130 & ~n1693;
  assign n1700 = pi005 & ~n1693;
  assign n1701 = pi005 & pi130;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1699 & n1702;
  assign n1704 = n1698 & n1703;
  assign n1705 = ~n1698 & ~n1703;
  assign n1706 = n1704 & ~n1705;
  assign n1707 = pi005 & ~n1706;
  assign n1708 = ~n355 & ~n1707;
  assign n1709 = pi012 & ~n1706;
  assign n1710 = n1708 & ~n1709;
  assign n1711 = n1685 & ~n1710;
  assign n1712 = ~n1684 & n1711;
  assign n1713 = pi005 & pi008;
  assign n1714 = ~n1700 & ~n1713;
  assign n1715 = ~n1694 & n1714;
  assign n1716 = ~pi005 & pi130;
  assign n1717 = ~n1695 & ~n1716;
  assign n1718 = ~n1699 & n1717;
  assign n1719 = ~n1715 & ~n1718;
  assign n1720 = ~n1673 & n1719;
  assign n1721 = ~n1683 & ~n1720;
  assign n1722 = ~n1681 & n1719;
  assign n1723 = n1721 & ~n1722;
  assign n1724 = ~n1719 & n1723;
  assign n1725 = n1719 & ~n1723;
  assign n1726 = n1724 & ~n1725;
  assign n1727 = ~n1684 & ~n1726;
  assign n1728 = ~n1712 & ~n1727;
  assign n1729 = n1711 & ~n1726;
  assign n1730 = n1728 & ~n1729;
  assign n1731 = ~n1684 & ~n1730;
  assign n1732 = ~n1656 & n1731;
  assign n1733 = ~n1665 & ~n1732;
  assign n1734 = ~n1664 & n1731;
  assign n1735 = n1733 & ~n1734;
  assign n1736 = ~n1648 & ~n1735;
  assign n1737 = n1656 & n1664;
  assign n1738 = ~n1665 & n1737;
  assign n1739 = ~n1706 & n1738;
  assign n1740 = n1637 & ~n1645;
  assign n1741 = ~n1637 & n1645;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = ~n1706 & ~n1742;
  assign n1744 = ~n1739 & ~n1743;
  assign n1745 = n1738 & ~n1742;
  assign n1746 = n1744 & ~n1745;
  assign n1747 = ~n1738 & ~n1746;
  assign n1748 = pi005 & pi048;
  assign n1749 = pi048 & n1748;
  assign n1750 = ~pi012 & pi031;
  assign n1751 = pi012 & ~pi031;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = pi048 & ~n1752;
  assign n1754 = ~n1749 & ~n1753;
  assign n1755 = n1748 & ~n1752;
  assign n1756 = n1754 & ~n1755;
  assign n1757 = ~n1747 & ~n1756;
  assign n1758 = ~n1684 & n1726;
  assign n1759 = ~n1656 & n1684;
  assign n1760 = ~n1665 & ~n1759;
  assign n1761 = ~n1664 & n1684;
  assign n1762 = n1760 & ~n1761;
  assign n1763 = n1758 & n1762;
  assign n1764 = ~n1756 & n1763;
  assign n1765 = ~n1757 & ~n1764;
  assign n1766 = ~n1747 & n1763;
  assign n1767 = n1765 & ~n1766;
  assign n1768 = n1747 & ~n1767;
  assign n1769 = ~n1637 & n1768;
  assign n1770 = ~n1647 & ~n1769;
  assign n1771 = ~n1645 & n1768;
  assign n1772 = n1770 & ~n1771;
  assign n1773 = ~n1768 & n1772;
  assign n1774 = n1768 & ~n1772;
  assign n1775 = n1773 & ~n1774;
  assign n1776 = n1736 & ~n1775;
  assign n1777 = n1628 & n1736;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = n1628 & ~n1775;
  assign n1780 = n1778 & ~n1779;
  assign n1781 = n1629 & ~n1780;
  assign n1782 = ~n1620 & n1781;
  assign n1783 = ~n1621 & ~n1782;
  assign n1784 = ~n1614 & n1781;
  assign n1785 = n1783 & ~n1784;
  assign n1786 = ~n1614 & n1785;
  assign n1787 = n1614 & ~n1785;
  assign n1788 = n1786 & ~n1787;
  assign n1789 = ~n1403 & ~n1788;
  assign n1790 = ~n1536 & ~n1789;
  assign n1791 = ~n1445 & n1453;
  assign n1792 = ~n1453 & n1791;
  assign n1793 = n1481 & n1489;
  assign n1794 = ~n1490 & n1793;
  assign n1795 = ~n1453 & ~n1794;
  assign n1796 = ~n1792 & ~n1795;
  assign n1797 = n1791 & ~n1794;
  assign n1798 = n1796 & ~n1797;
  assign n1799 = ~n1420 & ~n1798;
  assign n1800 = n1420 & ~n1506;
  assign n1801 = ~n1437 & ~n1523;
  assign n1802 = ~n1437 & ~n1497;
  assign n1803 = n1454 & ~n1497;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1437 & n1454;
  assign n1806 = n1804 & ~n1805;
  assign n1807 = n1801 & n1806;
  assign n1808 = n1420 & n1807;
  assign n1809 = ~n1800 & ~n1808;
  assign n1810 = ~n1506 & n1807;
  assign n1811 = n1809 & ~n1810;
  assign n1812 = n1799 & ~n1811;
  assign n1813 = ~n1788 & n1812;
  assign n1814 = n1789 & n1812;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1788 & n1789;
  assign n1817 = n1815 & ~n1816;
  assign n1818 = ~n1536 & ~n1817;
  assign n1819 = ~n1790 & ~n1818;
  assign n1820 = ~n1789 & ~n1817;
  assign n1821 = n1819 & ~n1820;
  assign n1822 = n1237 & ~n1245;
  assign n1823 = ~n1237 & n1245;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = n1220 & ~n1228;
  assign n1826 = ~n1220 & n1228;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = ~n1824 & ~n1827;
  assign n1829 = n1127 & n1828;
  assign n1830 = ~n1127 & n1277;
  assign n1831 = n1176 & ~n1195;
  assign n1832 = n1203 & ~n1211;
  assign n1833 = ~n1203 & n1211;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = n1176 & n1834;
  assign n1836 = ~n1831 & ~n1835;
  assign n1837 = ~n1195 & n1834;
  assign n1838 = n1836 & ~n1837;
  assign n1839 = ~n1195 & n1838;
  assign n1840 = ~n1167 & n1839;
  assign n1841 = n1167 & ~n1184;
  assign n1842 = n1167 & ~n1192;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = ~n1194 & n1843;
  assign n1845 = n1840 & n1844;
  assign n1846 = ~n1127 & n1845;
  assign n1847 = ~n1830 & ~n1846;
  assign n1848 = n1277 & n1845;
  assign n1849 = n1847 & ~n1848;
  assign n1850 = n1829 & ~n1849;
  assign n1851 = ~n1821 & n1850;
  assign n1852 = ~n1294 & ~n1821;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = ~n1294 & n1850;
  assign n1855 = n1853 & ~n1854;
  assign n1856 = n1294 & n1855;
  assign n1857 = ~n1294 & ~n1855;
  assign n1858 = n1856 & ~n1857;
  assign n1859 = ~n1063 & ~n1858;
  assign n1860 = pi058 & ~pi168;
  assign n1861 = ~pi005 & pi058;
  assign n1862 = pi005 & ~pi058;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = pi058 & ~n1863;
  assign n1865 = ~n1860 & ~n1864;
  assign n1866 = ~pi168 & ~n1863;
  assign n1867 = n1865 & ~n1866;
  assign n1868 = ~n381 & ~n1867;
  assign n1869 = n381 & n1867;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = pi005 & ~pi089;
  assign n1872 = ~n382 & ~n1871;
  assign n1873 = ~pi089 & n381;
  assign n1874 = n1872 & ~n1873;
  assign n1875 = ~n381 & n1874;
  assign n1876 = n381 & ~n1874;
  assign n1877 = n1875 & ~n1876;
  assign n1878 = pi047 & ~pi171;
  assign n1879 = ~pi005 & pi047;
  assign n1880 = pi005 & ~pi047;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = pi047 & ~n1881;
  assign n1883 = ~n1878 & ~n1882;
  assign n1884 = ~pi171 & ~n1881;
  assign n1885 = n1883 & ~n1884;
  assign n1886 = n1877 & ~n1885;
  assign n1887 = ~n1877 & n1885;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1870 & n1888;
  assign n1890 = ~n1870 & ~n1888;
  assign n1891 = n1889 & ~n1890;
  assign n1892 = ~n1063 & n1891;
  assign n1893 = ~n1859 & ~n1892;
  assign n1894 = ~n1858 & n1891;
  assign n1895 = n1893 & ~n1894;
  assign n1896 = n1063 & ~n1895;
  assign n1897 = ~pi174 & ~pi206;
  assign n1898 = pi174 & pi206;
  assign n1899 = n1897 & ~n1898;
  assign n1900 = pi011 & n1899;
  assign n1901 = pi166 & ~n1899;
  assign n1902 = ~n990 & ~n1901;
  assign n1903 = pi174 & ~n1899;
  assign n1904 = n1902 & ~n1903;
  assign n1905 = pi011 & ~n1904;
  assign n1906 = ~n1900 & ~n1905;
  assign n1907 = n1899 & ~n1904;
  assign n1908 = n1906 & ~n1907;
  assign n1909 = n1063 & ~n1868;
  assign n1910 = ~n1063 & n1868;
  assign n1911 = n1909 & ~n1910;
  assign n1912 = n1063 & ~n1911;
  assign n1913 = ~n381 & ~n1019;
  assign n1914 = ~pi005 & pi092;
  assign n1915 = ~pi005 & ~n1019;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = pi092 & ~n1019;
  assign n1918 = n1916 & ~n1917;
  assign n1919 = n1913 & ~n1918;
  assign n1920 = ~n1054 & n1919;
  assign n1921 = ~n1056 & n1919;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = ~n1054 & ~n1056;
  assign n1924 = n1922 & ~n1923;
  assign n1925 = n1054 & n1924;
  assign n1926 = ~n1054 & ~n1924;
  assign n1927 = n1925 & ~n1926;
  assign n1928 = ~n1011 & ~n1927;
  assign n1929 = n1063 & n1928;
  assign n1930 = ~n1912 & ~n1929;
  assign n1931 = ~n1911 & n1928;
  assign n1932 = n1930 & ~n1931;
  assign n1933 = n1877 & ~n1932;
  assign n1934 = ~n1886 & ~n1933;
  assign n1935 = ~n1885 & ~n1932;
  assign n1936 = n1934 & ~n1935;
  assign n1937 = n1908 & n1936;
  assign n1938 = ~n1908 & ~n1936;
  assign n1939 = n1937 & ~n1938;
  assign n1940 = n1896 & ~n1939;
  assign n1941 = ~n995 & n1896;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = ~n995 & ~n1939;
  assign n1944 = n1942 & ~n1943;
  assign po058 = ~n995 & ~n1944;
  assign n1946 = ~n786 & ~n834;
  assign n1947 = n797 & ~n846;
  assign n1948 = n797 & ~n831;
  assign n1949 = ~n797 & n831;
  assign n1950 = n1948 & ~n1949;
  assign n1951 = ~n846 & ~n1950;
  assign n1952 = ~n1947 & ~n1951;
  assign n1953 = n797 & ~n1950;
  assign n1954 = n1952 & ~n1953;
  assign n1955 = n1946 & ~n1954;
  assign n1956 = ~n1946 & n1954;
  assign po061 = ~n1955 & ~n1956;
  assign n1958 = ~n831 & n842;
  assign n1959 = n831 & ~n842;
  assign n1960 = n1958 & ~n1959;
  assign n1961 = n797 & ~n1960;
  assign n1962 = ~n797 & n1960;
  assign po062 = ~n1961 & ~n1962;
  assign n1964 = ~n821 & ~n828;
  assign n1965 = n821 & n828;
  assign n1966 = n1964 & ~n1965;
  assign n1967 = ~n835 & n1966;
  assign n1968 = n835 & ~n1966;
  assign n1969 = n1967 & ~n1968;
  assign n1970 = n811 & ~n1969;
  assign n1971 = ~n811 & n1969;
  assign po063 = ~n1970 & ~n1971;
  assign n1973 = pi205 & n360;
  assign n1974 = pi205 & n363;
  assign n1975 = pi205 & ~n1974;
  assign n1976 = ~n1973 & ~n1975;
  assign n1977 = n360 & ~n1974;
  assign n1978 = n1976 & ~n1977;
  assign n1979 = n823 & ~n1978;
  assign n1980 = ~n823 & n1978;
  assign po064 = ~n1979 & ~n1980;
  assign n1982 = n853 & n855;
  assign n1983 = ~n853 & ~n855;
  assign n1984 = n1982 & ~n1983;
  assign n1985 = ~n769 & ~n1984;
  assign n1986 = ~n855 & ~n857;
  assign n1987 = ~n855 & ~n1984;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = ~n857 & ~n1984;
  assign n1990 = n1988 & ~n1989;
  assign n1991 = ~n769 & n1990;
  assign n1992 = ~n1985 & ~n1991;
  assign n1993 = ~n1984 & n1990;
  assign n1994 = n1992 & ~n1993;
  assign n1995 = ~pi193 & ~n1994;
  assign n1996 = ~n742 & ~n1995;
  assign n1997 = ~n741 & ~n1994;
  assign n1998 = n1996 & ~n1997;
  assign n1999 = n733 & ~n1998;
  assign n2000 = ~n733 & n1998;
  assign po065 = ~n1999 & ~n2000;
  assign n2002 = n741 & ~n1994;
  assign n2003 = ~n741 & n1994;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = ~pi193 & ~n2004;
  assign n2006 = pi193 & n2004;
  assign po066 = ~n2005 & ~n2006;
  assign n2008 = ~pi191 & ~n853;
  assign n2009 = ~n765 & ~n2008;
  assign n2010 = ~n764 & ~n853;
  assign n2011 = n2009 & ~n2010;
  assign n2012 = n855 & ~n2011;
  assign n2013 = ~n855 & n2011;
  assign po067 = ~n2012 & ~n2013;
  assign n2015 = n853 & ~n857;
  assign n2016 = ~n853 & n857;
  assign po068 = ~n2015 & ~n2016;
  assign n2018 = ~n382 & ~n455;
  assign n2019 = pi132 & n381;
  assign n2020 = n2018 & ~n2019;
  assign n2021 = pi005 & n2020;
  assign n2022 = ~pi134 & pi135;
  assign n2023 = pi134 & ~pi135;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = pi005 & n2024;
  assign n2026 = ~n382 & ~n2025;
  assign n2027 = n381 & n2024;
  assign n2028 = n2026 & ~n2027;
  assign n2029 = pi005 & n2028;
  assign n2030 = ~pi136 & pi137;
  assign n2031 = pi136 & ~pi137;
  assign n2032 = ~n2030 & ~n2031;
  assign n2033 = pi005 & n2032;
  assign n2034 = ~n382 & ~n2033;
  assign n2035 = n381 & n2032;
  assign n2036 = n2034 & ~n2035;
  assign n2037 = pi005 & n2036;
  assign n2038 = ~pi138 & pi139;
  assign n2039 = pi138 & ~pi139;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = pi005 & n2040;
  assign n2042 = ~n382 & ~n2041;
  assign n2043 = n381 & n2040;
  assign n2044 = n2042 & ~n2043;
  assign n2045 = pi005 & n2044;
  assign n2046 = ~n2037 & n2045;
  assign n2047 = n2037 & ~n2045;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~n2029 & ~n2048;
  assign n2050 = n2029 & n2048;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = ~n2021 & ~n2051;
  assign n2053 = n2021 & n2051;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n607 & ~n902;
  assign n2056 = ~n607 & n902;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = n618 & ~n632;
  assign n2059 = ~n618 & n632;
  assign n2060 = ~n2058 & ~n2059;
  assign n2061 = n2057 & ~n2060;
  assign n2062 = ~n2057 & n2060;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = n687 & ~n2063;
  assign n2065 = ~n687 & n2063;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = pi060 & pi150;
  assign n2068 = ~pi005 & pi060;
  assign n2069 = pi005 & ~pi060;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = pi060 & ~n2070;
  assign n2072 = ~n2067 & ~n2071;
  assign n2073 = pi150 & ~n2070;
  assign n2074 = n2072 & ~n2073;
  assign n2075 = n669 & ~n2074;
  assign n2076 = ~n669 & n2074;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = n657 & ~n678;
  assign n2079 = ~n657 & n678;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = n2077 & ~n2080;
  assign n2082 = ~n2077 & n2080;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = n646 & ~n2083;
  assign n2085 = ~n646 & n2083;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = n2066 & ~n2086;
  assign n2088 = ~n2066 & n2086;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n2054 & ~n2089;
  assign n2091 = ~pi078 & pi079;
  assign n2092 = pi078 & ~pi079;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = pi005 & n2093;
  assign n2095 = ~n382 & ~n2094;
  assign n2096 = n381 & n2093;
  assign n2097 = n2095 & ~n2096;
  assign n2098 = pi005 & n2097;
  assign n2099 = pi070 & pi084;
  assign n2100 = ~pi005 & pi084;
  assign n2101 = pi005 & ~pi084;
  assign n2102 = ~n2100 & ~n2101;
  assign n2103 = pi070 & n2102;
  assign n2104 = ~n2099 & ~n2103;
  assign n2105 = pi084 & n2102;
  assign n2106 = n2104 & ~n2105;
  assign n2107 = n524 & ~n562;
  assign n2108 = ~n524 & n562;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = n2106 & ~n2109;
  assign n2111 = ~n2106 & n2109;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = ~pi076 & pi077;
  assign n2114 = pi076 & ~pi077;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = pi005 & n2115;
  assign n2117 = ~n382 & ~n2116;
  assign n2118 = n381 & n2115;
  assign n2119 = n2117 & ~n2118;
  assign n2120 = pi005 & n2119;
  assign n2121 = n551 & n2120;
  assign n2122 = ~n551 & ~n2120;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = n2112 & ~n2123;
  assign n2125 = ~n2112 & n2123;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n2098 & ~n2126;
  assign n2128 = n2098 & n2126;
  assign n2129 = ~n2127 & ~n2128;
  assign n2130 = n533 & ~n2129;
  assign n2131 = ~n533 & n2129;
  assign n2132 = ~n2130 & ~n2131;
  assign n2133 = n542 & ~n2132;
  assign n2134 = ~n542 & n2132;
  assign n2135 = ~n2133 & ~n2134;
  assign n2136 = ~n2089 & ~n2135;
  assign n2137 = ~n730 & n741;
  assign n2138 = n730 & ~n741;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = n755 & ~n2139;
  assign n2141 = ~n755 & n2139;
  assign n2142 = ~n2140 & ~n2141;
  assign n2143 = n764 & ~n2142;
  assign n2144 = ~n764 & n2142;
  assign n2145 = ~n2143 & ~n2144;
  assign n2146 = pi013 & pi162;
  assign n2147 = ~pi005 & pi013;
  assign n2148 = pi005 & ~pi013;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = pi013 & ~n2149;
  assign n2151 = ~n2146 & ~n2150;
  assign n2152 = pi162 & ~n2149;
  assign n2153 = n2151 & ~n2152;
  assign n2154 = n808 & ~n2153;
  assign n2155 = ~n808 & n2153;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = pi012 & pi152;
  assign n2158 = ~pi005 & pi012;
  assign n2159 = pi005 & ~pi012;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = pi012 & ~n2160;
  assign n2162 = ~n2157 & ~n2161;
  assign n2163 = pi152 & ~n2160;
  assign n2164 = n2162 & ~n2163;
  assign n2165 = n785 & ~n2164;
  assign n2166 = ~n785 & n2164;
  assign n2167 = ~n2165 & ~n2166;
  assign n2168 = n2156 & ~n2167;
  assign n2169 = ~n2156 & n2167;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = n820 & ~n2170;
  assign n2172 = ~n820 & n2170;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = n2145 & ~n2173;
  assign n2175 = ~n2145 & n2173;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = n794 & ~n2176;
  assign n2178 = ~n794 & n2176;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n2135 & n2179;
  assign n2181 = ~n2136 & ~n2180;
  assign n2182 = ~n2089 & n2179;
  assign n2183 = n2181 & ~n2182;
  assign po069 = ~n2090 | ~n2183;
  assign n2185 = n1329 & ~n1346;
  assign n2186 = ~n1329 & n1346;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = n1310 & ~n2187;
  assign n2189 = ~n1310 & n2187;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = n1360 & ~n2190;
  assign n2192 = ~n1360 & n2190;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = pi021 & ~pi195;
  assign n2195 = ~pi005 & pi021;
  assign n2196 = pi005 & ~pi021;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = pi021 & ~n2197;
  assign n2199 = ~n2194 & ~n2198;
  assign n2200 = ~pi195 & ~n2197;
  assign n2201 = n2199 & ~n2200;
  assign n2202 = n1453 & ~n2201;
  assign n2203 = ~n1453 & n2201;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = n2193 & ~n2204;
  assign n2206 = ~n2193 & n2204;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = n1463 & ~n2207;
  assign n2209 = ~n1463 & n2207;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = ~n1436 & n1489;
  assign n2212 = n1436 & ~n1489;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = n2210 & ~n2213;
  assign n2215 = ~n2210 & n2213;
  assign n2216 = ~n2214 & ~n2215;
  assign n2217 = n1419 & ~n2216;
  assign n2218 = ~n1419 & n2216;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = ~pi166 & pi174;
  assign n2221 = pi166 & ~pi174;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = ~pi005 & ~n2222;
  assign n2224 = pi005 & n2222;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = ~n2222 & ~n2225;
  assign n2227 = ~pi172 & pi173;
  assign n2228 = pi172 & ~pi173;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2222 & ~n2229;
  assign n2231 = ~n2226 & ~n2230;
  assign n2232 = ~n2225 & ~n2229;
  assign n2233 = n2231 & ~n2232;
  assign n2234 = pi059 & ~pi167;
  assign n2235 = ~pi005 & pi059;
  assign n2236 = pi005 & ~pi059;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = pi059 & ~n2237;
  assign n2239 = ~n2234 & ~n2238;
  assign n2240 = ~pi167 & ~n2237;
  assign n2241 = n2239 & ~n2240;
  assign n2242 = n1049 & ~n2241;
  assign n2243 = ~n1049 & n2241;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = n2233 & ~n2244;
  assign n2246 = ~n2233 & n2244;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = n1019 & ~n2247;
  assign n2249 = ~n1019 & n2247;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = n1010 & ~n1885;
  assign n2252 = ~n1010 & n1885;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = n2250 & ~n2253;
  assign n2255 = ~n2250 & n2253;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = n1867 & ~n2256;
  assign n2258 = ~n1867 & n2256;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = n1078 & ~n1142;
  assign n2261 = ~n1078 & n1142;
  assign n2262 = ~n2260 & ~n2261;
  assign n2263 = n1095 & ~n2262;
  assign n2264 = ~n1095 & n2262;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = n1111 & ~n2265;
  assign n2267 = ~n1111 & n2265;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = pi041 & ~pi175;
  assign n2270 = ~pi005 & pi041;
  assign n2271 = pi005 & ~pi041;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = pi041 & ~n2272;
  assign n2274 = ~n2269 & ~n2273;
  assign n2275 = ~pi175 & ~n2272;
  assign n2276 = n2274 & ~n2275;
  assign n2277 = pi027 & ~pi180;
  assign n2278 = pi005 & ~pi180;
  assign n2279 = ~n1150 & ~n2278;
  assign n2280 = pi027 & ~n2279;
  assign n2281 = ~n2277 & ~n2280;
  assign n2282 = ~pi180 & ~n2279;
  assign n2283 = n2281 & ~n2282;
  assign n2284 = n1245 & ~n2283;
  assign n2285 = ~n1245 & n2283;
  assign n2286 = ~n2284 & ~n2285;
  assign n2287 = n1192 & ~n2286;
  assign n2288 = ~n1192 & n2286;
  assign n2289 = ~n2287 & ~n2288;
  assign n2290 = n2276 & ~n2289;
  assign n2291 = ~n2276 & n2289;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = n1211 & ~n1228;
  assign n2294 = ~n1211 & n1228;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = n2292 & ~n2295;
  assign n2297 = ~n2292 & n2295;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = n2268 & ~n2298;
  assign n2300 = ~n2268 & n2298;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2259 & ~n2301;
  assign n2303 = n2219 & n2302;
  assign n2304 = pi031 & ~pi186;
  assign n2305 = pi005 & ~pi031;
  assign n2306 = ~n1685 & ~n2305;
  assign n2307 = pi031 & ~n2306;
  assign n2308 = ~n2304 & ~n2307;
  assign n2309 = ~pi186 & ~n2306;
  assign n2310 = n2308 & ~n2309;
  assign n2311 = n1681 & ~n1693;
  assign n2312 = ~n1681 & n1693;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = n2310 & ~n2313;
  assign n2315 = ~n2310 & n2313;
  assign n2316 = ~n2314 & ~n2315;
  assign n2317 = n1591 & ~n1608;
  assign n2318 = ~n1591 & n1608;
  assign n2319 = ~n2317 & ~n2318;
  assign n2320 = n1571 & ~n2319;
  assign n2321 = ~n1571 & n2319;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = n1552 & ~n2322;
  assign n2324 = ~n1552 & n2322;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = pi030 & ~pi185;
  assign n2327 = ~pi005 & pi030;
  assign n2328 = pi005 & ~pi030;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = pi030 & ~n2329;
  assign n2331 = ~n2326 & ~n2330;
  assign n2332 = ~pi185 & ~n2329;
  assign n2333 = n2331 & ~n2332;
  assign n2334 = n1645 & ~n2333;
  assign n2335 = ~n1645 & n2333;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = n2325 & ~n2336;
  assign n2338 = ~n2325 & n2336;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = n1664 & ~n2339;
  assign n2341 = ~n1664 & n2339;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = n2316 & ~n2342;
  assign n2344 = ~n2316 & n2342;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = n2302 & ~n2345;
  assign n2347 = ~n2303 & ~n2346;
  assign n2348 = n2219 & ~n2345;
  assign n2349 = n2347 & ~n2348;
  assign po070 = n2219 | n2349;
  assign n2351 = n1321 & ~n1338;
  assign n2352 = ~n1321 & n1338;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = n1302 & ~n2353;
  assign n2355 = ~n1302 & n2353;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = n1380 & ~n2356;
  assign n2358 = ~n1380 & n2356;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = pi050 & pi119;
  assign n2361 = pi005 & ~pi050;
  assign n2362 = ~n1498 & ~n2361;
  assign n2363 = pi050 & ~n2362;
  assign n2364 = ~n2360 & ~n2363;
  assign n2365 = pi119 & ~n2362;
  assign n2366 = n2364 & ~n2365;
  assign n2367 = n2359 & ~n2366;
  assign n2368 = ~n2359 & n2366;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = pi060 & pi120;
  assign n2371 = ~n2071 & ~n2370;
  assign n2372 = pi120 & ~n2070;
  assign n2373 = n2371 & ~n2372;
  assign n2374 = n1445 & ~n2373;
  assign n2375 = ~n1445 & n2373;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = ~n1428 & n1481;
  assign n2378 = n1428 & ~n1481;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = n2376 & ~n2379;
  assign n2381 = ~n2376 & n2379;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = n1411 & ~n2382;
  assign n2384 = ~n1411 & n2382;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = n2369 & n2385;
  assign n2387 = ~n2369 & ~n2385;
  assign n2388 = n2386 & ~n2387;
  assign n2389 = ~pi087 & pi088;
  assign n2390 = pi087 & ~pi088;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = pi005 & n2391;
  assign n2393 = ~n382 & ~n2392;
  assign n2394 = n381 & n2391;
  assign n2395 = n2393 & ~n2394;
  assign n2396 = pi005 & n2395;
  assign n2397 = ~pi089 & pi093;
  assign n2398 = pi089 & ~pi093;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = pi005 & ~n2399;
  assign n2401 = n996 & ~n2400;
  assign n2402 = ~n996 & n2400;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~n381 & ~n2403;
  assign n2405 = ~pi091 & pi092;
  assign n2406 = pi091 & ~pi092;
  assign n2407 = ~n2405 & ~n2406;
  assign n2408 = pi005 & n2407;
  assign n2409 = ~n382 & ~n2408;
  assign n2410 = n381 & n2407;
  assign n2411 = n2409 & ~n2410;
  assign n2412 = pi005 & n2411;
  assign n2413 = ~n2404 & n2412;
  assign n2414 = n2404 & ~n2412;
  assign n2415 = ~n2413 & ~n2414;
  assign n2416 = ~n2396 & ~n2415;
  assign n2417 = n2396 & n2415;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = ~n2369 & ~n2418;
  assign n2420 = ~n2385 & ~n2418;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = ~n2387 & n2421;
  assign n2423 = n2418 & n2422;
  assign n2424 = ~n2418 & ~n2422;
  assign n2425 = n2423 & ~n2424;
  assign n2426 = ~n2388 & ~n2425;
  assign n2427 = n1583 & ~n1600;
  assign n2428 = ~n1583 & n1600;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = n1563 & ~n2429;
  assign n2431 = ~n1563 & n2429;
  assign n2432 = ~n2430 & ~n2431;
  assign n2433 = n1544 & ~n2432;
  assign n2434 = ~n1544 & n2432;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = n1656 & ~n2435;
  assign n2437 = ~n1656 & n2435;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = pi013 & pi131;
  assign n2440 = ~n2150 & ~n2439;
  assign n2441 = pi131 & ~n2149;
  assign n2442 = n2440 & ~n2441;
  assign n2443 = n1673 & ~n2442;
  assign n2444 = ~n1673 & n2442;
  assign n2445 = ~n2443 & ~n2444;
  assign n2446 = pi008 & pi130;
  assign n2447 = pi005 & ~pi008;
  assign n2448 = ~n1696 & ~n2447;
  assign n2449 = pi008 & ~n2448;
  assign n2450 = ~n2446 & ~n2449;
  assign n2451 = pi130 & ~n2448;
  assign n2452 = n2450 & ~n2451;
  assign n2453 = n2445 & ~n2452;
  assign n2454 = ~n2445 & n2452;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = pi012 & pi121;
  assign n2457 = ~n2161 & ~n2456;
  assign n2458 = pi121 & ~n2160;
  assign n2459 = n2457 & ~n2458;
  assign n2460 = n1637 & ~n2459;
  assign n2461 = ~n1637 & n2459;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = n2455 & ~n2462;
  assign n2464 = ~n2455 & n2462;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = n2438 & ~n2465;
  assign n2467 = ~n2438 & n2465;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = ~n2388 & n2468;
  assign n2470 = ~n2426 & ~n2469;
  assign n2471 = ~n2425 & n2468;
  assign n2472 = n2470 & ~n2471;
  assign n2473 = ~n2388 & n2472;
  assign n2474 = ~pi098 & pi099;
  assign n2475 = pi098 & ~pi099;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = pi005 & n2476;
  assign n2478 = ~n382 & ~n2477;
  assign n2479 = n381 & n2476;
  assign n2480 = n2478 & ~n2479;
  assign n2481 = pi005 & n2480;
  assign n2482 = ~pi096 & pi097;
  assign n2483 = pi096 & ~pi097;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = pi005 & n2484;
  assign n2486 = ~n382 & ~n2485;
  assign n2487 = n381 & n2484;
  assign n2488 = n2486 & ~n2487;
  assign n2489 = pi005 & n2488;
  assign n2490 = ~n2481 & n2489;
  assign n2491 = n2481 & ~n2489;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = n1220 & ~n2492;
  assign n2494 = ~n1220 & n2492;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = pi070 & pi104;
  assign n2497 = ~pi005 & pi104;
  assign n2498 = pi005 & ~pi104;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = pi070 & n2499;
  assign n2501 = ~n2496 & ~n2500;
  assign n2502 = pi104 & n2499;
  assign n2503 = n2501 & ~n2502;
  assign n2504 = n1184 & ~n1237;
  assign n2505 = ~n1184 & n1237;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = n2503 & ~n2506;
  assign n2508 = ~n2503 & n2506;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = n1203 & ~n2509;
  assign n2511 = ~n1203 & n2509;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = n2495 & ~n2512;
  assign n2514 = ~n2495 & n2512;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n1157 & ~n2515;
  assign n2517 = ~n1157 & n2515;
  assign n2518 = ~n2516 & ~n2517;
  assign po071 = ~n2473 | ~n2518;
  assign n2520 = ~n925 & n935;
  assign n2521 = n925 & ~n935;
  assign po073 = ~n2520 & ~n2521;
  assign n2523 = ~n463 & ~n953;
  assign n2524 = n463 & n953;
  assign po074 = ~n2523 & ~n2524;
  assign n2526 = n1403 & n1813;
  assign n2527 = ~n1528 & ~n1813;
  assign n2528 = n1403 & n2527;
  assign n2529 = ~n2526 & ~n2528;
  assign n2530 = n1813 & n2527;
  assign n2531 = n2529 & ~n2530;
  assign n2532 = n1395 & n2531;
  assign n2533 = ~n1395 & ~n2531;
  assign po075 = ~n2532 | n2533;
  assign n2535 = ~n575 & ~n925;
  assign n2536 = ~n925 & ~n945;
  assign n2537 = ~n925 & ~n2536;
  assign n2538 = ~n2535 & ~n2537;
  assign n2539 = ~n575 & ~n2536;
  assign n2540 = n2538 & ~n2539;
  assign n2541 = n928 & ~n2540;
  assign n2542 = ~n928 & n2540;
  assign po077 = n2541 | n2542;
  assign n2544 = ~n554 & n935;
  assign n2545 = ~n554 & ~n925;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = ~n2520 & n2546;
  assign n2548 = n554 & ~n2547;
  assign n2549 = ~n571 & n2548;
  assign n2550 = ~n932 & n2548;
  assign n2551 = ~n571 & ~n2550;
  assign n2552 = ~n2549 & ~n2551;
  assign n2553 = n2548 & ~n2550;
  assign n2554 = n2552 & ~n2553;
  assign n2555 = n930 & ~n2554;
  assign n2556 = ~n930 & n2554;
  assign po078 = ~n2555 & ~n2556;
  assign n2558 = n567 & ~n2548;
  assign n2559 = ~n567 & n2548;
  assign n2560 = n2558 & ~n2559;
  assign n2561 = n932 & ~n2560;
  assign n2562 = ~n932 & n2560;
  assign po079 = ~n2561 & ~n2562;
  assign n2564 = ~pi176 & ~n925;
  assign n2565 = ~n563 & ~n2564;
  assign n2566 = ~n562 & ~n925;
  assign n2567 = n2565 & ~n2566;
  assign n2568 = n554 & ~n2567;
  assign n2569 = ~n554 & n2567;
  assign po080 = ~n2568 & ~n2569;
  assign n2571 = n453 & ~n963;
  assign n2572 = ~n436 & n453;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = ~n436 & ~n963;
  assign n2575 = n2573 & ~n2574;
  assign n2576 = ~n436 & ~n2575;
  assign n2577 = pi170 & n2576;
  assign n2578 = ~n444 & ~n2577;
  assign n2579 = ~n399 & n2576;
  assign n2580 = n2578 & ~n2579;
  assign n2581 = n469 & ~n953;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = n402 & n2581;
  assign n2584 = ~n2580 & n2583;
  assign n2585 = ~n2582 & ~n2584;
  assign n2586 = ~n2581 & n2583;
  assign n2587 = n2585 & ~n2586;
  assign n2588 = n392 & ~n2587;
  assign n2589 = ~n392 & n2587;
  assign po081 = ~n2588 & ~n2589;
  assign n2591 = n2576 & ~n2581;
  assign n2592 = n402 & n2591;
  assign n2593 = ~n402 & ~n2591;
  assign po082 = ~n2592 & ~n2593;
  assign n2595 = ~n421 & n953;
  assign n2596 = ~n2524 & ~n2595;
  assign n2597 = ~n421 & n463;
  assign n2598 = n2596 & ~n2597;
  assign n2599 = ~n421 & ~n2598;
  assign n2600 = pi169 & n2599;
  assign n2601 = ~n962 & ~n2600;
  assign n2602 = ~n428 & n2599;
  assign n2603 = n2601 & ~n2602;
  assign n2604 = n453 & ~n2603;
  assign n2605 = ~n453 & n2603;
  assign po083 = ~n2604 & ~n2605;
  assign n2607 = n431 & n2599;
  assign n2608 = ~n431 & ~n2599;
  assign po084 = ~n2607 & ~n2608;
  assign n2610 = ~po043 & ~po045;
  assign n2611 = ~po042 & po043;
  assign n2612 = ~po042 & ~po044;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = po043 & ~po044;
  assign n2615 = n2613 & ~n2614;
  assign n2616 = n2610 & ~n2615;
  assign n2617 = ~po070 & n2616;
  assign n2618 = ~po069 & po070;
  assign n2619 = ~po069 & ~po071;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = po070 & ~po071;
  assign n2622 = n2620 & ~n2621;
  assign po085 = ~n2617 | n2622;
  assign n2624 = ~n925 & n946;
  assign n2625 = n579 & n946;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = n579 & ~n925;
  assign n2628 = n2626 & ~n2627;
  assign n2629 = ~n579 & n2628;
  assign n2630 = n501 & ~n2629;
  assign n2631 = ~n590 & ~n2630;
  assign n2632 = pi183 & n2631;
  assign n2633 = ~n582 & ~n2632;
  assign n2634 = ~n477 & n2631;
  assign n2635 = n2633 & ~n2634;
  assign n2636 = n512 & ~n2635;
  assign n2637 = ~n512 & n2635;
  assign po087 = ~n2636 & ~n2637;
  assign n2639 = n480 & n2631;
  assign n2640 = ~n480 & ~n2631;
  assign po088 = ~n2639 & ~n2640;
  assign n2642 = pi181 & n2629;
  assign n2643 = ~n585 & ~n2642;
  assign n2644 = ~n497 & n2629;
  assign n2645 = n2643 & ~n2644;
  assign n2646 = n490 & ~n2645;
  assign n2647 = ~n490 & n2645;
  assign po089 = ~n2646 & ~n2647;
  assign n2649 = n497 & n2629;
  assign n2650 = ~n497 & ~n2629;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = ~pi181 & ~n2651;
  assign n2653 = pi181 & n2651;
  assign po090 = ~n2652 & ~n2653;
  assign n2655 = ~n711 & n873;
  assign n2656 = n711 & ~n873;
  assign po091 = ~n2655 & ~n2656;
  assign n2658 = ~pi011 & n974;
  assign n2659 = pi172 & pi206;
  assign n2660 = ~pi011 & n2659;
  assign n2661 = ~n2658 & ~n2660;
  assign n2662 = n974 & n2659;
  assign n2663 = n2661 & ~n2662;
  assign n2664 = pi173 & pi206;
  assign n2665 = n2663 & n2664;
  assign n2666 = ~n2663 & ~n2664;
  assign n2667 = ~n2665 & ~n2666;
  assign n2668 = ~pi011 & ~n2667;
  assign n2669 = pi011 & n2667;
  assign po092 = n2668 | n2669;
  assign n2671 = ~n974 & n2659;
  assign n2672 = n974 & ~n2659;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = ~pi011 & ~n2673;
  assign n2675 = pi011 & n2673;
  assign po094 = n2674 | n2675;
  assign n2677 = n688 & n709;
  assign n2678 = ~n695 & n709;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n688 & ~n695;
  assign n2681 = n2679 & ~n2680;
  assign n2682 = n695 & n2681;
  assign n2683 = ~n695 & ~n2681;
  assign n2684 = n2682 & ~n2683;
  assign n2685 = ~pi199 & ~n2684;
  assign n2686 = ~n658 & ~n2685;
  assign n2687 = ~n657 & ~n2684;
  assign n2688 = n2686 & ~n2687;
  assign n2689 = n719 & ~n873;
  assign n2690 = ~n2688 & n2689;
  assign n2691 = ~n660 & n2689;
  assign n2692 = ~n2688 & ~n2691;
  assign n2693 = ~n2690 & ~n2692;
  assign n2694 = n2689 & ~n2691;
  assign n2695 = n2693 & ~n2694;
  assign n2696 = n649 & ~n2695;
  assign n2697 = ~n649 & n2695;
  assign po096 = ~n2696 & ~n2697;
  assign n2699 = n2684 & ~n2689;
  assign n2700 = ~n2684 & n2689;
  assign n2701 = n2699 & ~n2700;
  assign n2702 = n660 & ~n2701;
  assign n2703 = ~n660 & n2701;
  assign po097 = ~n2702 & ~n2703;
  assign n2705 = ~pi196 & ~n873;
  assign n2706 = ~n679 & ~n2705;
  assign n2707 = ~n678 & ~n873;
  assign n2708 = n2706 & ~n2707;
  assign n2709 = ~pi197 & ~n2708;
  assign n2710 = ~n688 & ~n2709;
  assign n2711 = ~n687 & ~n2708;
  assign n2712 = n2710 & ~n2711;
  assign n2713 = n709 & ~n2712;
  assign n2714 = ~n709 & n2712;
  assign po098 = ~n2713 & ~n2714;
  assign n2716 = n690 & ~n2708;
  assign n2717 = ~n690 & n2708;
  assign po099 = ~n2716 & ~n2717;
  assign n2719 = n624 & ~n893;
  assign n2720 = n914 & ~n2719;
  assign n2721 = ~n914 & n2719;
  assign n2722 = n2720 & ~n2721;
  assign n2723 = ~pi203 & ~n2722;
  assign n2724 = ~n633 & ~n2723;
  assign n2725 = ~n632 & ~n2722;
  assign n2726 = n2724 & ~n2725;
  assign n2727 = n905 & ~n2726;
  assign n2728 = ~n905 & n2726;
  assign po100 = ~n2727 & ~n2728;
  assign n2730 = n635 & ~n2722;
  assign n2731 = ~n635 & n2722;
  assign po101 = ~n2730 & ~n2731;
  assign n2733 = ~pi201 & ~n893;
  assign n2734 = ~n619 & ~n2733;
  assign n2735 = ~n618 & ~n893;
  assign n2736 = n2734 & ~n2735;
  assign n2737 = n610 & ~n2736;
  assign n2738 = ~n610 & n2736;
  assign po102 = ~n2737 & ~n2738;
  assign n2740 = ~n618 & n893;
  assign n2741 = n618 & ~n893;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = ~pi201 & ~n2742;
  assign n2744 = pi201 & n2742;
  assign po103 = ~n2743 & ~n2744;
  assign n2746 = n590 & ~n594;
  assign n2747 = ~n590 & n594;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = n512 & ~n2748;
  assign n2750 = ~n512 & n2748;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = n585 & n2751;
  assign n2753 = ~n585 & ~n2751;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = n490 & ~n2754;
  assign n2756 = ~n490 & n2754;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = ~n501 & ~n590;
  assign n2759 = ~pi183 & n2758;
  assign n2760 = ~n478 & ~n2759;
  assign n2761 = ~n477 & n2758;
  assign n2762 = n2760 & ~n2761;
  assign n2763 = n477 & ~n2762;
  assign n2764 = ~n477 & n2762;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = n512 & ~n2765;
  assign n2767 = ~n512 & n2765;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = n586 & ~n2768;
  assign n2770 = ~n586 & n2768;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = n490 & ~n2771;
  assign n2773 = ~n490 & n2771;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = n2757 & ~n2774;
  assign n2776 = ~n2629 & ~n2774;
  assign n2777 = n2629 & n2774;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = n2757 & ~n2778;
  assign n2780 = ~n2775 & ~n2779;
  assign n2781 = ~n2774 & ~n2778;
  assign n2782 = n2780 & ~n2781;
  assign n2783 = n480 & ~n2782;
  assign n2784 = ~n480 & n2782;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = pi177 & n563;
  assign n2787 = ~n553 & ~n2786;
  assign n2788 = n551 & n563;
  assign n2789 = n2787 & ~n2788;
  assign n2790 = n575 & ~n2789;
  assign n2791 = ~n575 & n2789;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = ~pi178 & n552;
  assign n2794 = ~n543 & ~n2793;
  assign n2795 = ~n542 & n552;
  assign n2796 = n2794 & ~n2795;
  assign n2797 = ~n563 & ~n2796;
  assign n2798 = n935 & n2797;
  assign n2799 = ~n935 & ~n2797;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = n563 & n571;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = n930 & n2802;
  assign n2804 = ~n930 & ~n2802;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = n932 & ~n2805;
  assign n2807 = ~n932 & n2805;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = n2792 & ~n2808;
  assign n2810 = ~n2792 & n2808;
  assign n2811 = ~n2809 & ~n2810;
  assign n2812 = n928 & ~n2811;
  assign n2813 = ~n928 & n2811;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = n571 & ~n942;
  assign n2816 = pi179 & n2815;
  assign n2817 = ~n929 & ~n2816;
  assign n2818 = n533 & n2815;
  assign n2819 = n2817 & ~n2818;
  assign n2820 = ~n2815 & ~n2819;
  assign n2821 = n2815 & n2819;
  assign n2822 = ~n2820 & ~n2821;
  assign n2823 = pi177 & n934;
  assign n2824 = ~n553 & ~n2823;
  assign n2825 = n551 & n934;
  assign n2826 = n2824 & ~n2825;
  assign n2827 = ~n554 & ~n563;
  assign n2828 = ~n564 & ~n2827;
  assign n2829 = n930 & ~n2828;
  assign n2830 = ~n930 & n2828;
  assign n2831 = ~n2829 & ~n2830;
  assign n2832 = n932 & ~n2831;
  assign n2833 = ~n932 & n2831;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = n2826 & ~n2834;
  assign n2836 = ~n2826 & n2834;
  assign n2837 = ~n2835 & ~n2836;
  assign n2838 = n2822 & ~n2837;
  assign n2839 = ~n2822 & n2837;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = n928 & ~n2840;
  assign n2842 = ~n928 & n2840;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = ~n2814 & n2843;
  assign n2845 = n925 & ~n2843;
  assign n2846 = ~n925 & n2843;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = ~n2814 & ~n2847;
  assign n2849 = ~n2844 & ~n2848;
  assign n2850 = n2843 & ~n2847;
  assign n2851 = n2849 & ~n2850;
  assign n2852 = n2785 & ~n2851;
  assign n2853 = ~n2785 & n2851;
  assign po104 = ~n2852 & ~n2853;
  assign n2855 = pi011 & ~pi206;
  assign n2856 = ~n989 & ~n2855;
  assign n2857 = pi011 & ~n2856;
  assign n2858 = pi172 & n2856;
  assign n2859 = ~n2659 & ~n2858;
  assign n2860 = pi206 & n2856;
  assign n2861 = n2859 & ~n2860;
  assign n2862 = ~pi173 & ~n2861;
  assign n2863 = pi173 & n2861;
  assign n2864 = ~n2862 & ~n2863;
  assign n2865 = pi011 & ~n2864;
  assign n2866 = ~n2857 & ~n2865;
  assign n2867 = ~n2856 & ~n2864;
  assign n2868 = n2866 & ~n2867;
  assign n2869 = n2664 & ~n2868;
  assign n2870 = pi011 & ~n2659;
  assign n2871 = ~n2660 & ~n2870;
  assign n2872 = ~n974 & ~n2871;
  assign n2873 = ~n2868 & ~n2872;
  assign n2874 = n2868 & n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = n2664 & ~n2875;
  assign n2877 = ~n2869 & ~n2876;
  assign n2878 = ~n2868 & ~n2875;
  assign n2879 = n2877 & ~n2878;
  assign n2880 = pi053 & ~n963;
  assign n2881 = ~n411 & ~n2880;
  assign n2882 = ~n410 & ~n963;
  assign n2883 = n2881 & ~n2882;
  assign n2884 = ~n421 & ~n2883;
  assign n2885 = n463 & n2884;
  assign n2886 = ~n463 & ~n2884;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = ~n421 & n2887;
  assign n2889 = ~n2576 & ~n2884;
  assign n2890 = n2576 & n2884;
  assign n2891 = n2889 & ~n2890;
  assign n2892 = ~n421 & ~n2891;
  assign n2893 = ~n2888 & ~n2892;
  assign n2894 = n2887 & ~n2891;
  assign n2895 = n2893 & ~n2894;
  assign n2896 = n2887 & ~n2895;
  assign n2897 = pi169 & n421;
  assign n2898 = ~n962 & ~n2897;
  assign n2899 = n421 & ~n428;
  assign n2900 = n2898 & ~n2899;
  assign n2901 = n2580 & ~n2900;
  assign n2902 = ~n2580 & n2900;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = ~n402 & n453;
  assign n2905 = ~n967 & ~n2904;
  assign n2906 = n2903 & ~n2905;
  assign n2907 = ~n2903 & n2905;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = n392 & ~n2908;
  assign n2910 = ~n392 & n2908;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = ~n2896 & ~n2911;
  assign n2913 = n2896 & n2911;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = n431 & ~n453;
  assign n2916 = ~n467 & ~n2915;
  assign n2917 = n421 & ~n2916;
  assign n2918 = ~n421 & n2916;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = ~n469 & n2576;
  assign n2921 = pi170 & ~n2920;
  assign n2922 = ~n444 & ~n2921;
  assign n2923 = ~n399 & ~n2920;
  assign n2924 = n2922 & ~n2923;
  assign n2925 = ~n2920 & ~n2924;
  assign n2926 = n2920 & n2924;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = pi169 & n2597;
  assign n2929 = ~n962 & ~n2928;
  assign n2930 = ~n428 & n2597;
  assign n2931 = n2929 & ~n2930;
  assign n2932 = n392 & ~n2931;
  assign n2933 = ~n392 & n2931;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = n2927 & ~n2934;
  assign n2936 = ~n2927 & n2934;
  assign n2937 = ~n2935 & ~n2936;
  assign n2938 = n2919 & ~n2937;
  assign n2939 = ~n2919 & n2937;
  assign n2940 = ~n2938 & ~n2939;
  assign n2941 = n2914 & ~n2940;
  assign n2942 = ~n953 & ~n2940;
  assign n2943 = n953 & n2940;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = n2914 & ~n2944;
  assign n2946 = ~n2941 & ~n2945;
  assign n2947 = ~n2940 & ~n2944;
  assign n2948 = n2946 & ~n2947;
  assign n2949 = n2879 & ~n2948;
  assign n2950 = ~n2879 & n2948;
  assign po105 = n2949 | n2950;
  assign n2952 = pi203 & ~n632;
  assign n2953 = pi203 & ~n914;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = ~n917 & n2954;
  assign n2956 = n632 & ~n2955;
  assign n2957 = ~n632 & n2955;
  assign n2958 = ~n2956 & ~n2957;
  assign n2959 = n905 & ~n2958;
  assign n2960 = ~n905 & n2958;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = n620 & n2961;
  assign n2963 = ~n620 & ~n2961;
  assign n2964 = ~n2962 & ~n2963;
  assign n2965 = n610 & ~n2964;
  assign n2966 = ~n610 & n2964;
  assign n2967 = ~n2965 & ~n2966;
  assign n2968 = ~n624 & n914;
  assign n2969 = pi203 & n2968;
  assign n2970 = ~n2952 & ~n2969;
  assign n2971 = ~n632 & n2968;
  assign n2972 = n2970 & ~n2971;
  assign n2973 = ~pi203 & ~n2972;
  assign n2974 = pi203 & n2972;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = n905 & ~n2975;
  assign n2977 = ~n905 & n2975;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = ~n619 & ~n2978;
  assign n2980 = n619 & n2978;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = n610 & ~n2981;
  assign n2983 = ~n610 & n2981;
  assign n2984 = ~n2982 & ~n2983;
  assign n2985 = ~n2967 & ~n2984;
  assign n2986 = n893 & ~n2984;
  assign n2987 = ~n893 & n2984;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = ~n2967 & n2988;
  assign n2990 = ~n2985 & ~n2989;
  assign n2991 = ~n2984 & n2988;
  assign n2992 = n2990 & ~n2991;
  assign n2993 = n635 & ~n2992;
  assign n2994 = ~n635 & n2992;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = n678 & ~n2684;
  assign n2997 = ~pi198 & n688;
  assign n2998 = ~n670 & ~n2997;
  assign n2999 = ~n669 & n688;
  assign n3000 = n2998 & ~n2999;
  assign n3001 = ~n679 & n3000;
  assign n3002 = n679 & ~n3000;
  assign n3003 = n3001 & ~n3002;
  assign n3004 = n678 & ~n3003;
  assign n3005 = ~n2996 & ~n3004;
  assign n3006 = ~n2684 & ~n3003;
  assign n3007 = n3005 & ~n3006;
  assign n3008 = ~n678 & ~n3007;
  assign n3009 = ~n678 & n3003;
  assign n3010 = ~n3004 & ~n3009;
  assign n3011 = ~pi196 & ~n3010;
  assign n3012 = pi196 & n3010;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = ~n3008 & n3013;
  assign n3015 = n3008 & ~n3013;
  assign n3016 = n3014 & ~n3015;
  assign n3017 = pi197 & n679;
  assign n3018 = ~n689 & ~n3017;
  assign n3019 = n679 & n687;
  assign n3020 = n3018 & ~n3019;
  assign n3021 = n2688 & ~n3020;
  assign n3022 = ~n2688 & n3020;
  assign n3023 = ~n3021 & ~n3022;
  assign n3024 = n3016 & ~n3023;
  assign n3025 = ~n3016 & n3023;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = n649 & ~n3026;
  assign n3028 = ~n649 & n3026;
  assign n3029 = ~n3027 & ~n3028;
  assign n3030 = n660 & ~n3029;
  assign n3031 = ~n660 & n3029;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = n709 & ~n3032;
  assign n3034 = ~n709 & n3032;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = n873 & ~n3035;
  assign n3037 = pi197 & n710;
  assign n3038 = ~n689 & ~n3037;
  assign n3039 = n687 & n710;
  assign n3040 = n3038 & ~n3039;
  assign n3041 = ~n719 & n2684;
  assign n3042 = pi199 & n3041;
  assign n3043 = ~n659 & ~n3042;
  assign n3044 = n657 & n3041;
  assign n3045 = n3043 & ~n3044;
  assign n3046 = ~n3041 & ~n3045;
  assign n3047 = n3041 & n3045;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = n649 & ~n3048;
  assign n3050 = ~n649 & n3048;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = n3040 & ~n3051;
  assign n3053 = ~n3040 & n3051;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = n690 & ~n709;
  assign n3056 = ~n715 & ~n3055;
  assign n3057 = n660 & ~n3056;
  assign n3058 = ~n660 & n3056;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n679 & ~n3059;
  assign n3061 = n679 & n3059;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n3054 & ~n3062;
  assign n3064 = ~n3054 & n3062;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = ~n873 & n3065;
  assign n3067 = ~n3036 & ~n3066;
  assign n3068 = n3036 & n3066;
  assign n3069 = n3067 & ~n3068;
  assign n3070 = n2995 & ~n3069;
  assign n3071 = ~n2995 & n3069;
  assign po106 = n3070 | n3071;
  assign n3073 = pi193 & ~n741;
  assign n3074 = pi193 & n769;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = ~n741 & n769;
  assign n3077 = n3075 & ~n3076;
  assign n3078 = n741 & ~n3077;
  assign n3079 = ~n741 & n3077;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = n733 & ~n3080;
  assign n3082 = ~n733 & n3080;
  assign n3083 = ~n3081 & ~n3082;
  assign n3084 = n855 & ~n3083;
  assign n3085 = ~n855 & n3083;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = ~n856 & ~n3086;
  assign n3088 = n856 & n3086;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = n853 & ~n3089;
  assign n3091 = ~n733 & n741;
  assign n3092 = n733 & ~n741;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = ~pi193 & ~n3093;
  assign n3095 = pi193 & n3093;
  assign n3096 = ~n3094 & ~n3095;
  assign n3097 = ~n765 & ~n3096;
  assign n3098 = n765 & n3096;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = n855 & ~n3099;
  assign n3101 = ~n855 & n3099;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = pi192 & n856;
  assign n3104 = ~n854 & ~n3103;
  assign n3105 = n755 & n856;
  assign n3106 = n3104 & ~n3105;
  assign n3107 = pi193 & ~n3106;
  assign n3108 = ~n743 & ~n3107;
  assign n3109 = n741 & ~n3106;
  assign n3110 = n3108 & ~n3109;
  assign n3111 = n3106 & ~n3110;
  assign n3112 = ~n3106 & n3110;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = n3102 & ~n3113;
  assign n3115 = ~n3102 & n3113;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = ~n853 & ~n3116;
  assign n3118 = ~n3090 & ~n3117;
  assign n3119 = n3090 & n3117;
  assign n3120 = n3118 & ~n3119;
  assign n3121 = n811 & ~n3120;
  assign n3122 = ~n811 & n3120;
  assign n3123 = ~n3121 & ~n3122;
  assign n3124 = n797 & ~n3123;
  assign n3125 = ~n797 & n3123;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = ~n360 & n363;
  assign n3128 = ~pi187 & n3127;
  assign n3129 = ~n821 & ~n3128;
  assign n3130 = ~n820 & n3127;
  assign n3131 = n3129 & ~n3130;
  assign n3132 = n795 & n846;
  assign n3133 = ~n366 & n823;
  assign n3134 = ~n366 & ~n811;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = ~n811 & n823;
  assign n3137 = n3135 & ~n3136;
  assign n3138 = n823 & n3137;
  assign n3139 = ~n823 & ~n3137;
  assign n3140 = n3138 & ~n3139;
  assign n3141 = ~n795 & ~n3140;
  assign n3142 = n795 & n3141;
  assign n3143 = ~n3132 & ~n3142;
  assign n3144 = n846 & n3141;
  assign n3145 = n3143 & ~n3144;
  assign n3146 = n1946 & ~n3145;
  assign n3147 = ~n1946 & n3145;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = ~n363 & ~n842;
  assign n3150 = n363 & n842;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = n842 & ~n3151;
  assign n3153 = n363 & ~n3140;
  assign n3154 = n363 & n3151;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n3140 & n3151;
  assign n3157 = n3155 & ~n3156;
  assign n3158 = ~n360 & ~n3157;
  assign n3159 = n360 & n3157;
  assign n3160 = ~n3158 & ~n3159;
  assign n3161 = n842 & ~n3160;
  assign n3162 = ~n3152 & ~n3161;
  assign n3163 = ~n3151 & ~n3160;
  assign n3164 = n3162 & ~n3163;
  assign n3165 = n3148 & ~n3164;
  assign n3166 = ~n3148 & n3164;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = n3131 & ~n3167;
  assign n3169 = ~n3131 & n3167;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = n360 & ~n842;
  assign n3172 = ~n360 & n3171;
  assign n3173 = ~pi188 & n821;
  assign n3174 = ~n809 & ~n3173;
  assign n3175 = ~n808 & n821;
  assign n3176 = n3174 & ~n3175;
  assign n3177 = ~n360 & ~n3176;
  assign n3178 = n366 & n3177;
  assign n3179 = ~n366 & ~n3177;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = ~n360 & ~n3180;
  assign n3182 = ~n3172 & ~n3181;
  assign n3183 = n3171 & ~n3180;
  assign n3184 = n3182 & ~n3183;
  assign n3185 = pi187 & n360;
  assign n3186 = ~n822 & ~n3185;
  assign n3187 = n360 & n820;
  assign n3188 = n3186 & ~n3187;
  assign n3189 = n3184 & ~n3188;
  assign n3190 = ~n3184 & n3188;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = n846 & ~n3191;
  assign n3193 = ~n846 & n3191;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = n1946 & ~n3194;
  assign n3196 = ~n1946 & n3194;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = n3170 & ~n3197;
  assign n3199 = ~pi205 & ~n3197;
  assign n3200 = pi205 & n3197;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = n3170 & ~n3201;
  assign n3203 = ~n3198 & ~n3202;
  assign n3204 = ~n3197 & ~n3201;
  assign n3205 = n3203 & ~n3204;
  assign n3206 = n3126 & ~n3205;
  assign n3207 = ~n3126 & n3205;
  assign po107 = n3206 | n3207;
  assign po037 = ~pi004;
  assign po000 = pi164;
  assign po001 = pi000;
  assign po002 = pi000;
  assign po003 = pi167;
  assign po004 = pi169;
  assign po005 = pi170;
  assign po006 = pi171;
  assign po007 = pi172;
  assign po008 = pi173;
  assign po009 = pi175;
  assign po010 = pi177;
  assign po011 = pi178;
  assign po012 = pi179;
  assign po013 = pi180;
  assign po014 = pi181;
  assign po015 = pi182;
  assign po016 = pi183;
  assign po017 = pi184;
  assign po018 = pi185;
  assign po019 = pi186;
  assign po020 = pi187;
  assign po021 = pi188;
  assign po022 = pi189;
  assign po023 = pi190;
  assign po024 = pi191;
  assign po025 = pi192;
  assign po026 = pi193;
  assign po027 = pi194;
  assign po028 = pi195;
  assign po029 = pi197;
  assign po030 = pi198;
  assign po031 = pi199;
  assign po032 = pi200;
  assign po033 = pi201;
  assign po034 = pi202;
  assign po035 = pi203;
  assign po036 = pi204;
  assign po038 = pi168;
  assign po039 = pi176;
  assign po040 = pi196;
  assign po046 = pi000;
  assign po047 = pi053;
  assign po049 = po037;
  assign po050 = po048;
  assign po052 = po037;
  assign po053 = po051;
  assign po054 = pi000;
  assign po059 = po058;
  assign po060 = po057;
  assign po072 = po058;
  assign po076 = po057;
  assign po086 = po057;
  assign po093 = po092;
  assign po095 = po094;
endmodule


