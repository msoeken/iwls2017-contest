// Benchmark "mesh10" written by ABC on Wed Apr 26 18:30:59 2017

module mesh10 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    po0  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419;
  output po0;
  wire n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
  assign n422 = pi409 & pi419;
  assign n423 = pi398 & n422;
  assign n424 = ~pi398 & pi419;
  assign n425 = ~n423 & ~n424;
  assign n426 = pi399 & n425;
  assign n427 = ~pi399 & ~n425;
  assign n428 = ~n426 & ~n427;
  assign n429 = pi408 & ~n428;
  assign n430 = pi358 & n429;
  assign n431 = ~pi358 & ~n428;
  assign n432 = ~n430 & ~n431;
  assign n433 = pi359 & n432;
  assign n434 = ~pi359 & ~n432;
  assign n435 = ~n433 & ~n434;
  assign n436 = pi407 & ~n435;
  assign n437 = pi318 & n436;
  assign n438 = ~pi318 & ~n435;
  assign n439 = ~n437 & ~n438;
  assign n440 = pi319 & n439;
  assign n441 = ~pi319 & ~n439;
  assign n442 = ~n440 & ~n441;
  assign n443 = pi406 & ~n442;
  assign n444 = pi278 & n443;
  assign n445 = ~pi278 & ~n442;
  assign n446 = ~n444 & ~n445;
  assign n447 = pi279 & n446;
  assign n448 = ~pi279 & ~n446;
  assign n449 = ~n447 & ~n448;
  assign n450 = pi405 & ~n449;
  assign n451 = pi238 & n450;
  assign n452 = ~pi238 & ~n449;
  assign n453 = ~n451 & ~n452;
  assign n454 = pi239 & n453;
  assign n455 = ~pi239 & ~n453;
  assign n456 = ~n454 & ~n455;
  assign n457 = pi404 & ~n456;
  assign n458 = pi198 & n457;
  assign n459 = ~pi198 & ~n456;
  assign n460 = ~n458 & ~n459;
  assign n461 = pi199 & n460;
  assign n462 = ~pi199 & ~n460;
  assign n463 = ~n461 & ~n462;
  assign n464 = pi403 & ~n463;
  assign n465 = pi158 & n464;
  assign n466 = ~pi158 & ~n463;
  assign n467 = ~n465 & ~n466;
  assign n468 = pi159 & n467;
  assign n469 = ~pi159 & ~n467;
  assign n470 = ~n468 & ~n469;
  assign n471 = pi402 & ~n470;
  assign n472 = pi118 & n471;
  assign n473 = ~pi118 & ~n470;
  assign n474 = ~n472 & ~n473;
  assign n475 = pi119 & n474;
  assign n476 = ~pi119 & ~n474;
  assign n477 = ~n475 & ~n476;
  assign n478 = pi401 & ~n477;
  assign n479 = pi078 & n478;
  assign n480 = ~pi078 & ~n477;
  assign n481 = ~n479 & ~n480;
  assign n482 = pi079 & n481;
  assign n483 = ~pi079 & ~n481;
  assign n484 = ~n482 & ~n483;
  assign n485 = pi036 & pi400;
  assign n486 = ~n484 & n485;
  assign n487 = ~pi036 & pi400;
  assign n488 = ~n486 & ~n487;
  assign n489 = pi037 & n488;
  assign n490 = ~pi037 & ~n488;
  assign n491 = ~n489 & ~n490;
  assign n492 = pi076 & n478;
  assign n493 = ~pi076 & pi401;
  assign n494 = ~n492 & ~n493;
  assign n495 = pi077 & n494;
  assign n496 = ~pi077 & ~n494;
  assign n497 = ~n495 & ~n496;
  assign n498 = pi116 & n471;
  assign n499 = ~pi116 & pi402;
  assign n500 = ~n498 & ~n499;
  assign n501 = pi117 & n500;
  assign n502 = ~pi117 & ~n500;
  assign n503 = ~n501 & ~n502;
  assign n504 = pi156 & n464;
  assign n505 = ~pi156 & pi403;
  assign n506 = ~n504 & ~n505;
  assign n507 = pi157 & n506;
  assign n508 = ~pi157 & ~n506;
  assign n509 = ~n507 & ~n508;
  assign n510 = pi196 & n457;
  assign n511 = ~pi196 & pi404;
  assign n512 = ~n510 & ~n511;
  assign n513 = pi197 & n512;
  assign n514 = ~pi197 & ~n512;
  assign n515 = ~n513 & ~n514;
  assign n516 = pi236 & n450;
  assign n517 = ~pi236 & pi405;
  assign n518 = ~n516 & ~n517;
  assign n519 = pi237 & n518;
  assign n520 = ~pi237 & ~n518;
  assign n521 = ~n519 & ~n520;
  assign n522 = pi276 & n443;
  assign n523 = ~pi276 & pi406;
  assign n524 = ~n522 & ~n523;
  assign n525 = pi277 & n524;
  assign n526 = ~pi277 & ~n524;
  assign n527 = ~n525 & ~n526;
  assign n528 = pi316 & n436;
  assign n529 = ~pi316 & pi407;
  assign n530 = ~n528 & ~n529;
  assign n531 = pi317 & n530;
  assign n532 = ~pi317 & ~n530;
  assign n533 = ~n531 & ~n532;
  assign n534 = pi356 & n429;
  assign n535 = ~pi356 & pi408;
  assign n536 = ~n534 & ~n535;
  assign n537 = pi357 & n536;
  assign n538 = ~pi357 & ~n536;
  assign n539 = ~n537 & ~n538;
  assign n540 = pi396 & n422;
  assign n541 = ~pi396 & pi409;
  assign n542 = ~n540 & ~n541;
  assign n543 = pi397 & n542;
  assign n544 = ~pi397 & ~n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = pi418 & ~n545;
  assign n547 = pi394 & n546;
  assign n548 = ~pi394 & pi418;
  assign n549 = ~n547 & ~n548;
  assign n550 = pi395 & n549;
  assign n551 = ~pi395 & ~n549;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n539 & ~n552;
  assign n554 = pi354 & n553;
  assign n555 = ~pi354 & ~n552;
  assign n556 = ~n554 & ~n555;
  assign n557 = pi355 & n556;
  assign n558 = ~pi355 & ~n556;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n533 & ~n559;
  assign n561 = pi314 & n560;
  assign n562 = ~pi314 & ~n559;
  assign n563 = ~n561 & ~n562;
  assign n564 = pi315 & n563;
  assign n565 = ~pi315 & ~n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n527 & ~n566;
  assign n568 = pi274 & n567;
  assign n569 = ~pi274 & ~n566;
  assign n570 = ~n568 & ~n569;
  assign n571 = pi275 & n570;
  assign n572 = ~pi275 & ~n570;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n521 & ~n573;
  assign n575 = pi234 & n574;
  assign n576 = ~pi234 & ~n573;
  assign n577 = ~n575 & ~n576;
  assign n578 = pi235 & n577;
  assign n579 = ~pi235 & ~n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n515 & ~n580;
  assign n582 = pi194 & n581;
  assign n583 = ~pi194 & ~n580;
  assign n584 = ~n582 & ~n583;
  assign n585 = pi195 & n584;
  assign n586 = ~pi195 & ~n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n509 & ~n587;
  assign n589 = pi154 & n588;
  assign n590 = ~pi154 & ~n587;
  assign n591 = ~n589 & ~n590;
  assign n592 = pi155 & n591;
  assign n593 = ~pi155 & ~n591;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n503 & ~n594;
  assign n596 = pi114 & n595;
  assign n597 = ~pi114 & ~n594;
  assign n598 = ~n596 & ~n597;
  assign n599 = pi115 & n598;
  assign n600 = ~pi115 & ~n598;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n497 & ~n601;
  assign n603 = pi074 & n602;
  assign n604 = ~pi074 & ~n601;
  assign n605 = ~n603 & ~n604;
  assign n606 = pi075 & n605;
  assign n607 = ~pi075 & ~n605;
  assign n608 = ~n606 & ~n607;
  assign n609 = pi032 & ~n491;
  assign n610 = ~n608 & n609;
  assign n611 = ~pi032 & ~n491;
  assign n612 = ~n610 & ~n611;
  assign n613 = pi033 & n612;
  assign n614 = ~pi033 & ~n612;
  assign n615 = ~n613 & ~n614;
  assign n616 = pi072 & n602;
  assign n617 = ~pi072 & ~n497;
  assign n618 = ~n616 & ~n617;
  assign n619 = pi073 & n618;
  assign n620 = ~pi073 & ~n618;
  assign n621 = ~n619 & ~n620;
  assign n622 = pi112 & n595;
  assign n623 = ~pi112 & ~n503;
  assign n624 = ~n622 & ~n623;
  assign n625 = pi113 & n624;
  assign n626 = ~pi113 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = pi152 & n588;
  assign n629 = ~pi152 & ~n509;
  assign n630 = ~n628 & ~n629;
  assign n631 = pi153 & n630;
  assign n632 = ~pi153 & ~n630;
  assign n633 = ~n631 & ~n632;
  assign n634 = pi192 & n581;
  assign n635 = ~pi192 & ~n515;
  assign n636 = ~n634 & ~n635;
  assign n637 = pi193 & n636;
  assign n638 = ~pi193 & ~n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = pi232 & n574;
  assign n641 = ~pi232 & ~n521;
  assign n642 = ~n640 & ~n641;
  assign n643 = pi233 & n642;
  assign n644 = ~pi233 & ~n642;
  assign n645 = ~n643 & ~n644;
  assign n646 = pi272 & n567;
  assign n647 = ~pi272 & ~n527;
  assign n648 = ~n646 & ~n647;
  assign n649 = pi273 & n648;
  assign n650 = ~pi273 & ~n648;
  assign n651 = ~n649 & ~n650;
  assign n652 = pi312 & n560;
  assign n653 = ~pi312 & ~n533;
  assign n654 = ~n652 & ~n653;
  assign n655 = pi313 & n654;
  assign n656 = ~pi313 & ~n654;
  assign n657 = ~n655 & ~n656;
  assign n658 = pi352 & n553;
  assign n659 = ~pi352 & ~n539;
  assign n660 = ~n658 & ~n659;
  assign n661 = pi353 & n660;
  assign n662 = ~pi353 & ~n660;
  assign n663 = ~n661 & ~n662;
  assign n664 = pi392 & n546;
  assign n665 = ~pi392 & ~n545;
  assign n666 = ~n664 & ~n665;
  assign n667 = pi393 & n666;
  assign n668 = ~pi393 & ~n666;
  assign n669 = ~n667 & ~n668;
  assign n670 = pi417 & ~n669;
  assign n671 = pi390 & n670;
  assign n672 = ~pi390 & pi417;
  assign n673 = ~n671 & ~n672;
  assign n674 = pi391 & n673;
  assign n675 = ~pi391 & ~n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n663 & ~n676;
  assign n678 = pi350 & n677;
  assign n679 = ~pi350 & ~n676;
  assign n680 = ~n678 & ~n679;
  assign n681 = pi351 & n680;
  assign n682 = ~pi351 & ~n680;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n657 & ~n683;
  assign n685 = pi310 & n684;
  assign n686 = ~pi310 & ~n683;
  assign n687 = ~n685 & ~n686;
  assign n688 = pi311 & n687;
  assign n689 = ~pi311 & ~n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n651 & ~n690;
  assign n692 = pi270 & n691;
  assign n693 = ~pi270 & ~n690;
  assign n694 = ~n692 & ~n693;
  assign n695 = pi271 & n694;
  assign n696 = ~pi271 & ~n694;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n645 & ~n697;
  assign n699 = pi230 & n698;
  assign n700 = ~pi230 & ~n697;
  assign n701 = ~n699 & ~n700;
  assign n702 = pi231 & n701;
  assign n703 = ~pi231 & ~n701;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~n639 & ~n704;
  assign n706 = pi190 & n705;
  assign n707 = ~pi190 & ~n704;
  assign n708 = ~n706 & ~n707;
  assign n709 = pi191 & n708;
  assign n710 = ~pi191 & ~n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n633 & ~n711;
  assign n713 = pi150 & n712;
  assign n714 = ~pi150 & ~n711;
  assign n715 = ~n713 & ~n714;
  assign n716 = pi151 & n715;
  assign n717 = ~pi151 & ~n715;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n627 & ~n718;
  assign n720 = pi110 & n719;
  assign n721 = ~pi110 & ~n718;
  assign n722 = ~n720 & ~n721;
  assign n723 = pi111 & n722;
  assign n724 = ~pi111 & ~n722;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n621 & ~n725;
  assign n727 = pi070 & n726;
  assign n728 = ~pi070 & ~n725;
  assign n729 = ~n727 & ~n728;
  assign n730 = pi071 & n729;
  assign n731 = ~pi071 & ~n729;
  assign n732 = ~n730 & ~n731;
  assign n733 = pi028 & ~n615;
  assign n734 = ~n732 & n733;
  assign n735 = ~pi028 & ~n615;
  assign n736 = ~n734 & ~n735;
  assign n737 = pi029 & n736;
  assign n738 = ~pi029 & ~n736;
  assign n739 = ~n737 & ~n738;
  assign n740 = pi068 & n726;
  assign n741 = ~pi068 & ~n621;
  assign n742 = ~n740 & ~n741;
  assign n743 = pi069 & n742;
  assign n744 = ~pi069 & ~n742;
  assign n745 = ~n743 & ~n744;
  assign n746 = pi108 & n719;
  assign n747 = ~pi108 & ~n627;
  assign n748 = ~n746 & ~n747;
  assign n749 = pi109 & n748;
  assign n750 = ~pi109 & ~n748;
  assign n751 = ~n749 & ~n750;
  assign n752 = pi148 & n712;
  assign n753 = ~pi148 & ~n633;
  assign n754 = ~n752 & ~n753;
  assign n755 = pi149 & n754;
  assign n756 = ~pi149 & ~n754;
  assign n757 = ~n755 & ~n756;
  assign n758 = pi188 & n705;
  assign n759 = ~pi188 & ~n639;
  assign n760 = ~n758 & ~n759;
  assign n761 = pi189 & n760;
  assign n762 = ~pi189 & ~n760;
  assign n763 = ~n761 & ~n762;
  assign n764 = pi228 & n698;
  assign n765 = ~pi228 & ~n645;
  assign n766 = ~n764 & ~n765;
  assign n767 = pi229 & n766;
  assign n768 = ~pi229 & ~n766;
  assign n769 = ~n767 & ~n768;
  assign n770 = pi268 & n691;
  assign n771 = ~pi268 & ~n651;
  assign n772 = ~n770 & ~n771;
  assign n773 = pi269 & n772;
  assign n774 = ~pi269 & ~n772;
  assign n775 = ~n773 & ~n774;
  assign n776 = pi308 & n684;
  assign n777 = ~pi308 & ~n657;
  assign n778 = ~n776 & ~n777;
  assign n779 = pi309 & n778;
  assign n780 = ~pi309 & ~n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = pi348 & n677;
  assign n783 = ~pi348 & ~n663;
  assign n784 = ~n782 & ~n783;
  assign n785 = pi349 & n784;
  assign n786 = ~pi349 & ~n784;
  assign n787 = ~n785 & ~n786;
  assign n788 = pi388 & n670;
  assign n789 = ~pi388 & ~n669;
  assign n790 = ~n788 & ~n789;
  assign n791 = pi389 & n790;
  assign n792 = ~pi389 & ~n790;
  assign n793 = ~n791 & ~n792;
  assign n794 = pi416 & ~n793;
  assign n795 = pi386 & n794;
  assign n796 = ~pi386 & pi416;
  assign n797 = ~n795 & ~n796;
  assign n798 = pi387 & n797;
  assign n799 = ~pi387 & ~n797;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~n787 & ~n800;
  assign n802 = pi346 & n801;
  assign n803 = ~pi346 & ~n800;
  assign n804 = ~n802 & ~n803;
  assign n805 = pi347 & n804;
  assign n806 = ~pi347 & ~n804;
  assign n807 = ~n805 & ~n806;
  assign n808 = ~n781 & ~n807;
  assign n809 = pi306 & n808;
  assign n810 = ~pi306 & ~n807;
  assign n811 = ~n809 & ~n810;
  assign n812 = pi307 & n811;
  assign n813 = ~pi307 & ~n811;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n775 & ~n814;
  assign n816 = pi266 & n815;
  assign n817 = ~pi266 & ~n814;
  assign n818 = ~n816 & ~n817;
  assign n819 = pi267 & n818;
  assign n820 = ~pi267 & ~n818;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~n769 & ~n821;
  assign n823 = pi226 & n822;
  assign n824 = ~pi226 & ~n821;
  assign n825 = ~n823 & ~n824;
  assign n826 = pi227 & n825;
  assign n827 = ~pi227 & ~n825;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n763 & ~n828;
  assign n830 = pi186 & n829;
  assign n831 = ~pi186 & ~n828;
  assign n832 = ~n830 & ~n831;
  assign n833 = pi187 & n832;
  assign n834 = ~pi187 & ~n832;
  assign n835 = ~n833 & ~n834;
  assign n836 = ~n757 & ~n835;
  assign n837 = pi146 & n836;
  assign n838 = ~pi146 & ~n835;
  assign n839 = ~n837 & ~n838;
  assign n840 = pi147 & n839;
  assign n841 = ~pi147 & ~n839;
  assign n842 = ~n840 & ~n841;
  assign n843 = ~n751 & ~n842;
  assign n844 = pi106 & n843;
  assign n845 = ~pi106 & ~n842;
  assign n846 = ~n844 & ~n845;
  assign n847 = pi107 & n846;
  assign n848 = ~pi107 & ~n846;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~n745 & ~n849;
  assign n851 = pi066 & n850;
  assign n852 = ~pi066 & ~n849;
  assign n853 = ~n851 & ~n852;
  assign n854 = pi067 & n853;
  assign n855 = ~pi067 & ~n853;
  assign n856 = ~n854 & ~n855;
  assign n857 = pi024 & ~n739;
  assign n858 = ~n856 & n857;
  assign n859 = ~pi024 & ~n739;
  assign n860 = ~n858 & ~n859;
  assign n861 = pi025 & n860;
  assign n862 = ~pi025 & ~n860;
  assign n863 = ~n861 & ~n862;
  assign n864 = pi064 & n850;
  assign n865 = ~pi064 & ~n745;
  assign n866 = ~n864 & ~n865;
  assign n867 = pi065 & n866;
  assign n868 = ~pi065 & ~n866;
  assign n869 = ~n867 & ~n868;
  assign n870 = pi104 & n843;
  assign n871 = ~pi104 & ~n751;
  assign n872 = ~n870 & ~n871;
  assign n873 = pi105 & n872;
  assign n874 = ~pi105 & ~n872;
  assign n875 = ~n873 & ~n874;
  assign n876 = pi144 & n836;
  assign n877 = ~pi144 & ~n757;
  assign n878 = ~n876 & ~n877;
  assign n879 = pi145 & n878;
  assign n880 = ~pi145 & ~n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = pi184 & n829;
  assign n883 = ~pi184 & ~n763;
  assign n884 = ~n882 & ~n883;
  assign n885 = pi185 & n884;
  assign n886 = ~pi185 & ~n884;
  assign n887 = ~n885 & ~n886;
  assign n888 = pi224 & n822;
  assign n889 = ~pi224 & ~n769;
  assign n890 = ~n888 & ~n889;
  assign n891 = pi225 & n890;
  assign n892 = ~pi225 & ~n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = pi264 & n815;
  assign n895 = ~pi264 & ~n775;
  assign n896 = ~n894 & ~n895;
  assign n897 = pi265 & n896;
  assign n898 = ~pi265 & ~n896;
  assign n899 = ~n897 & ~n898;
  assign n900 = pi304 & n808;
  assign n901 = ~pi304 & ~n781;
  assign n902 = ~n900 & ~n901;
  assign n903 = pi305 & n902;
  assign n904 = ~pi305 & ~n902;
  assign n905 = ~n903 & ~n904;
  assign n906 = pi344 & n801;
  assign n907 = ~pi344 & ~n787;
  assign n908 = ~n906 & ~n907;
  assign n909 = pi345 & n908;
  assign n910 = ~pi345 & ~n908;
  assign n911 = ~n909 & ~n910;
  assign n912 = pi384 & n794;
  assign n913 = ~pi384 & ~n793;
  assign n914 = ~n912 & ~n913;
  assign n915 = pi385 & n914;
  assign n916 = ~pi385 & ~n914;
  assign n917 = ~n915 & ~n916;
  assign n918 = pi415 & ~n917;
  assign n919 = pi382 & n918;
  assign n920 = ~pi382 & pi415;
  assign n921 = ~n919 & ~n920;
  assign n922 = pi383 & n921;
  assign n923 = ~pi383 & ~n921;
  assign n924 = ~n922 & ~n923;
  assign n925 = ~n911 & ~n924;
  assign n926 = pi342 & n925;
  assign n927 = ~pi342 & ~n924;
  assign n928 = ~n926 & ~n927;
  assign n929 = pi343 & n928;
  assign n930 = ~pi343 & ~n928;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n905 & ~n931;
  assign n933 = pi302 & n932;
  assign n934 = ~pi302 & ~n931;
  assign n935 = ~n933 & ~n934;
  assign n936 = pi303 & n935;
  assign n937 = ~pi303 & ~n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n899 & ~n938;
  assign n940 = pi262 & n939;
  assign n941 = ~pi262 & ~n938;
  assign n942 = ~n940 & ~n941;
  assign n943 = pi263 & n942;
  assign n944 = ~pi263 & ~n942;
  assign n945 = ~n943 & ~n944;
  assign n946 = ~n893 & ~n945;
  assign n947 = pi222 & n946;
  assign n948 = ~pi222 & ~n945;
  assign n949 = ~n947 & ~n948;
  assign n950 = pi223 & n949;
  assign n951 = ~pi223 & ~n949;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n887 & ~n952;
  assign n954 = pi182 & n953;
  assign n955 = ~pi182 & ~n952;
  assign n956 = ~n954 & ~n955;
  assign n957 = pi183 & n956;
  assign n958 = ~pi183 & ~n956;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n881 & ~n959;
  assign n961 = pi142 & n960;
  assign n962 = ~pi142 & ~n959;
  assign n963 = ~n961 & ~n962;
  assign n964 = pi143 & n963;
  assign n965 = ~pi143 & ~n963;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n875 & ~n966;
  assign n968 = pi102 & n967;
  assign n969 = ~pi102 & ~n966;
  assign n970 = ~n968 & ~n969;
  assign n971 = pi103 & n970;
  assign n972 = ~pi103 & ~n970;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n869 & ~n973;
  assign n975 = pi062 & n974;
  assign n976 = ~pi062 & ~n973;
  assign n977 = ~n975 & ~n976;
  assign n978 = pi063 & n977;
  assign n979 = ~pi063 & ~n977;
  assign n980 = ~n978 & ~n979;
  assign n981 = pi020 & ~n863;
  assign n982 = ~n980 & n981;
  assign n983 = ~pi020 & ~n863;
  assign n984 = ~n982 & ~n983;
  assign n985 = pi021 & n984;
  assign n986 = ~pi021 & ~n984;
  assign n987 = ~n985 & ~n986;
  assign n988 = pi060 & n974;
  assign n989 = ~pi060 & ~n869;
  assign n990 = ~n988 & ~n989;
  assign n991 = pi061 & n990;
  assign n992 = ~pi061 & ~n990;
  assign n993 = ~n991 & ~n992;
  assign n994 = pi100 & n967;
  assign n995 = ~pi100 & ~n875;
  assign n996 = ~n994 & ~n995;
  assign n997 = pi101 & n996;
  assign n998 = ~pi101 & ~n996;
  assign n999 = ~n997 & ~n998;
  assign n1000 = pi140 & n960;
  assign n1001 = ~pi140 & ~n881;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = pi141 & n1002;
  assign n1004 = ~pi141 & ~n1002;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = pi180 & n953;
  assign n1007 = ~pi180 & ~n887;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = pi181 & n1008;
  assign n1010 = ~pi181 & ~n1008;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = pi220 & n946;
  assign n1013 = ~pi220 & ~n893;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = pi221 & n1014;
  assign n1016 = ~pi221 & ~n1014;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = pi260 & n939;
  assign n1019 = ~pi260 & ~n899;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = pi261 & n1020;
  assign n1022 = ~pi261 & ~n1020;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = pi300 & n932;
  assign n1025 = ~pi300 & ~n905;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = pi301 & n1026;
  assign n1028 = ~pi301 & ~n1026;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = pi340 & n925;
  assign n1031 = ~pi340 & ~n911;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = pi341 & n1032;
  assign n1034 = ~pi341 & ~n1032;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = pi380 & n918;
  assign n1037 = ~pi380 & ~n917;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = pi381 & n1038;
  assign n1040 = ~pi381 & ~n1038;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = pi414 & ~n1041;
  assign n1043 = pi378 & n1042;
  assign n1044 = ~pi378 & pi414;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = pi379 & n1045;
  assign n1047 = ~pi379 & ~n1045;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1035 & ~n1048;
  assign n1050 = pi338 & n1049;
  assign n1051 = ~pi338 & ~n1048;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = pi339 & n1052;
  assign n1054 = ~pi339 & ~n1052;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1029 & ~n1055;
  assign n1057 = pi298 & n1056;
  assign n1058 = ~pi298 & ~n1055;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = pi299 & n1059;
  assign n1061 = ~pi299 & ~n1059;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1023 & ~n1062;
  assign n1064 = pi258 & n1063;
  assign n1065 = ~pi258 & ~n1062;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = pi259 & n1066;
  assign n1068 = ~pi259 & ~n1066;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = ~n1017 & ~n1069;
  assign n1071 = pi218 & n1070;
  assign n1072 = ~pi218 & ~n1069;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = pi219 & n1073;
  assign n1075 = ~pi219 & ~n1073;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = ~n1011 & ~n1076;
  assign n1078 = pi178 & n1077;
  assign n1079 = ~pi178 & ~n1076;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = pi179 & n1080;
  assign n1082 = ~pi179 & ~n1080;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n1005 & ~n1083;
  assign n1085 = pi138 & n1084;
  assign n1086 = ~pi138 & ~n1083;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = pi139 & n1087;
  assign n1089 = ~pi139 & ~n1087;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = ~n999 & ~n1090;
  assign n1092 = pi098 & n1091;
  assign n1093 = ~pi098 & ~n1090;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = pi099 & n1094;
  assign n1096 = ~pi099 & ~n1094;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = ~n993 & ~n1097;
  assign n1099 = pi058 & n1098;
  assign n1100 = ~pi058 & ~n1097;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = pi059 & n1101;
  assign n1103 = ~pi059 & ~n1101;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = pi016 & ~n987;
  assign n1106 = ~n1104 & n1105;
  assign n1107 = ~pi016 & ~n987;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = pi017 & n1108;
  assign n1110 = ~pi017 & ~n1108;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = pi056 & n1098;
  assign n1113 = ~pi056 & ~n993;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = pi057 & n1114;
  assign n1116 = ~pi057 & ~n1114;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = pi096 & n1091;
  assign n1119 = ~pi096 & ~n999;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = pi097 & n1120;
  assign n1122 = ~pi097 & ~n1120;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = pi136 & n1084;
  assign n1125 = ~pi136 & ~n1005;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = pi137 & n1126;
  assign n1128 = ~pi137 & ~n1126;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = pi176 & n1077;
  assign n1131 = ~pi176 & ~n1011;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = pi177 & n1132;
  assign n1134 = ~pi177 & ~n1132;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = pi216 & n1070;
  assign n1137 = ~pi216 & ~n1017;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = pi217 & n1138;
  assign n1140 = ~pi217 & ~n1138;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = pi256 & n1063;
  assign n1143 = ~pi256 & ~n1023;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = pi257 & n1144;
  assign n1146 = ~pi257 & ~n1144;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = pi296 & n1056;
  assign n1149 = ~pi296 & ~n1029;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = pi297 & n1150;
  assign n1152 = ~pi297 & ~n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = pi336 & n1049;
  assign n1155 = ~pi336 & ~n1035;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = pi337 & n1156;
  assign n1158 = ~pi337 & ~n1156;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = pi376 & n1042;
  assign n1161 = ~pi376 & ~n1041;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = pi377 & n1162;
  assign n1164 = ~pi377 & ~n1162;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = pi413 & ~n1165;
  assign n1167 = pi374 & n1166;
  assign n1168 = ~pi374 & pi413;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = pi375 & n1169;
  assign n1171 = ~pi375 & ~n1169;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n1159 & ~n1172;
  assign n1174 = pi334 & n1173;
  assign n1175 = ~pi334 & ~n1172;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = pi335 & n1176;
  assign n1178 = ~pi335 & ~n1176;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = ~n1153 & ~n1179;
  assign n1181 = pi294 & n1180;
  assign n1182 = ~pi294 & ~n1179;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = pi295 & n1183;
  assign n1185 = ~pi295 & ~n1183;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = ~n1147 & ~n1186;
  assign n1188 = pi254 & n1187;
  assign n1189 = ~pi254 & ~n1186;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = pi255 & n1190;
  assign n1192 = ~pi255 & ~n1190;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1141 & ~n1193;
  assign n1195 = pi214 & n1194;
  assign n1196 = ~pi214 & ~n1193;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = pi215 & n1197;
  assign n1199 = ~pi215 & ~n1197;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1135 & ~n1200;
  assign n1202 = pi174 & n1201;
  assign n1203 = ~pi174 & ~n1200;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = pi175 & n1204;
  assign n1206 = ~pi175 & ~n1204;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~n1129 & ~n1207;
  assign n1209 = pi134 & n1208;
  assign n1210 = ~pi134 & ~n1207;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = pi135 & n1211;
  assign n1213 = ~pi135 & ~n1211;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1123 & ~n1214;
  assign n1216 = pi094 & n1215;
  assign n1217 = ~pi094 & ~n1214;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = pi095 & n1218;
  assign n1220 = ~pi095 & ~n1218;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n1117 & ~n1221;
  assign n1223 = pi054 & n1222;
  assign n1224 = ~pi054 & ~n1221;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = pi055 & n1225;
  assign n1227 = ~pi055 & ~n1225;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = pi012 & ~n1111;
  assign n1230 = ~n1228 & n1229;
  assign n1231 = ~pi012 & ~n1111;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = pi013 & n1232;
  assign n1234 = ~pi013 & ~n1232;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = pi052 & n1222;
  assign n1237 = ~pi052 & ~n1117;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = pi053 & n1238;
  assign n1240 = ~pi053 & ~n1238;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = pi092 & n1215;
  assign n1243 = ~pi092 & ~n1123;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = pi093 & n1244;
  assign n1246 = ~pi093 & ~n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = pi132 & n1208;
  assign n1249 = ~pi132 & ~n1129;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = pi133 & n1250;
  assign n1252 = ~pi133 & ~n1250;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = pi172 & n1201;
  assign n1255 = ~pi172 & ~n1135;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = pi173 & n1256;
  assign n1258 = ~pi173 & ~n1256;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = pi212 & n1194;
  assign n1261 = ~pi212 & ~n1141;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = pi213 & n1262;
  assign n1264 = ~pi213 & ~n1262;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = pi252 & n1187;
  assign n1267 = ~pi252 & ~n1147;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = pi253 & n1268;
  assign n1270 = ~pi253 & ~n1268;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = pi292 & n1180;
  assign n1273 = ~pi292 & ~n1153;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = pi293 & n1274;
  assign n1276 = ~pi293 & ~n1274;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = pi332 & n1173;
  assign n1279 = ~pi332 & ~n1159;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = pi333 & n1280;
  assign n1282 = ~pi333 & ~n1280;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = pi372 & n1166;
  assign n1285 = ~pi372 & ~n1165;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = pi373 & n1286;
  assign n1288 = ~pi373 & ~n1286;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = pi412 & ~n1289;
  assign n1291 = pi370 & n1290;
  assign n1292 = ~pi370 & pi412;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = pi371 & n1293;
  assign n1295 = ~pi371 & ~n1293;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~n1283 & ~n1296;
  assign n1298 = pi330 & n1297;
  assign n1299 = ~pi330 & ~n1296;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = pi331 & n1300;
  assign n1302 = ~pi331 & ~n1300;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~n1277 & ~n1303;
  assign n1305 = pi290 & n1304;
  assign n1306 = ~pi290 & ~n1303;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = pi291 & n1307;
  assign n1309 = ~pi291 & ~n1307;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1271 & ~n1310;
  assign n1312 = pi250 & n1311;
  assign n1313 = ~pi250 & ~n1310;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = pi251 & n1314;
  assign n1316 = ~pi251 & ~n1314;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = ~n1265 & ~n1317;
  assign n1319 = pi210 & n1318;
  assign n1320 = ~pi210 & ~n1317;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = pi211 & n1321;
  assign n1323 = ~pi211 & ~n1321;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n1259 & ~n1324;
  assign n1326 = pi170 & n1325;
  assign n1327 = ~pi170 & ~n1324;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = pi171 & n1328;
  assign n1330 = ~pi171 & ~n1328;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = ~n1253 & ~n1331;
  assign n1333 = pi130 & n1332;
  assign n1334 = ~pi130 & ~n1331;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = pi131 & n1335;
  assign n1337 = ~pi131 & ~n1335;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~n1247 & ~n1338;
  assign n1340 = pi090 & n1339;
  assign n1341 = ~pi090 & ~n1338;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = pi091 & n1342;
  assign n1344 = ~pi091 & ~n1342;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1241 & ~n1345;
  assign n1347 = pi050 & n1346;
  assign n1348 = ~pi050 & ~n1345;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = pi051 & n1349;
  assign n1351 = ~pi051 & ~n1349;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = pi008 & ~n1235;
  assign n1354 = ~n1352 & n1353;
  assign n1355 = ~pi008 & ~n1235;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = pi009 & n1356;
  assign n1358 = ~pi009 & ~n1356;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = pi048 & n1346;
  assign n1361 = ~pi048 & ~n1241;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = pi049 & n1362;
  assign n1364 = ~pi049 & ~n1362;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = pi088 & n1339;
  assign n1367 = ~pi088 & ~n1247;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = pi089 & n1368;
  assign n1370 = ~pi089 & ~n1368;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = pi128 & n1332;
  assign n1373 = ~pi128 & ~n1253;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = pi129 & n1374;
  assign n1376 = ~pi129 & ~n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = pi168 & n1325;
  assign n1379 = ~pi168 & ~n1259;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = pi169 & n1380;
  assign n1382 = ~pi169 & ~n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = pi208 & n1318;
  assign n1385 = ~pi208 & ~n1265;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = pi209 & n1386;
  assign n1388 = ~pi209 & ~n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = pi248 & n1311;
  assign n1391 = ~pi248 & ~n1271;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = pi249 & n1392;
  assign n1394 = ~pi249 & ~n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = pi288 & n1304;
  assign n1397 = ~pi288 & ~n1277;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = pi289 & n1398;
  assign n1400 = ~pi289 & ~n1398;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = pi328 & n1297;
  assign n1403 = ~pi328 & ~n1283;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = pi329 & n1404;
  assign n1406 = ~pi329 & ~n1404;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = pi368 & n1290;
  assign n1409 = ~pi368 & ~n1289;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = pi369 & n1410;
  assign n1412 = ~pi369 & ~n1410;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = pi411 & ~n1413;
  assign n1415 = pi366 & n1414;
  assign n1416 = ~pi366 & pi411;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = pi367 & n1417;
  assign n1419 = ~pi367 & ~n1417;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = ~n1407 & ~n1420;
  assign n1422 = pi326 & n1421;
  assign n1423 = ~pi326 & ~n1420;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = pi327 & n1424;
  assign n1426 = ~pi327 & ~n1424;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1401 & ~n1427;
  assign n1429 = pi286 & n1428;
  assign n1430 = ~pi286 & ~n1427;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = pi287 & n1431;
  assign n1433 = ~pi287 & ~n1431;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n1395 & ~n1434;
  assign n1436 = pi246 & n1435;
  assign n1437 = ~pi246 & ~n1434;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = pi247 & n1438;
  assign n1440 = ~pi247 & ~n1438;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~n1389 & ~n1441;
  assign n1443 = pi206 & n1442;
  assign n1444 = ~pi206 & ~n1441;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = pi207 & n1445;
  assign n1447 = ~pi207 & ~n1445;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1383 & ~n1448;
  assign n1450 = pi166 & n1449;
  assign n1451 = ~pi166 & ~n1448;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = pi167 & n1452;
  assign n1454 = ~pi167 & ~n1452;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~n1377 & ~n1455;
  assign n1457 = pi126 & n1456;
  assign n1458 = ~pi126 & ~n1455;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = pi127 & n1459;
  assign n1461 = ~pi127 & ~n1459;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = ~n1371 & ~n1462;
  assign n1464 = pi086 & n1463;
  assign n1465 = ~pi086 & ~n1462;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = pi087 & n1466;
  assign n1468 = ~pi087 & ~n1466;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = ~n1365 & ~n1469;
  assign n1471 = pi046 & n1470;
  assign n1472 = ~pi046 & ~n1469;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = pi047 & n1473;
  assign n1475 = ~pi047 & ~n1473;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = pi004 & ~n1359;
  assign n1478 = ~n1476 & n1477;
  assign n1479 = ~pi004 & ~n1359;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = pi005 & n1480;
  assign n1482 = ~pi005 & ~n1480;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = pi044 & n1470;
  assign n1485 = ~pi044 & ~n1365;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = pi045 & n1486;
  assign n1488 = ~pi045 & ~n1486;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = pi084 & n1463;
  assign n1491 = ~pi084 & ~n1371;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = pi085 & n1492;
  assign n1494 = ~pi085 & ~n1492;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = pi124 & n1456;
  assign n1497 = ~pi124 & ~n1377;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = pi125 & n1498;
  assign n1500 = ~pi125 & ~n1498;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = pi164 & n1449;
  assign n1503 = ~pi164 & ~n1383;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = pi165 & n1504;
  assign n1506 = ~pi165 & ~n1504;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = pi204 & n1442;
  assign n1509 = ~pi204 & ~n1389;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = pi205 & n1510;
  assign n1512 = ~pi205 & ~n1510;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = pi244 & n1435;
  assign n1515 = ~pi244 & ~n1395;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = pi245 & n1516;
  assign n1518 = ~pi245 & ~n1516;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = pi284 & n1428;
  assign n1521 = ~pi284 & ~n1401;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = pi285 & n1522;
  assign n1524 = ~pi285 & ~n1522;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = pi324 & n1421;
  assign n1527 = ~pi324 & ~n1407;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = pi325 & n1528;
  assign n1530 = ~pi325 & ~n1528;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = pi364 & n1414;
  assign n1533 = ~pi364 & ~n1413;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = pi365 & n1534;
  assign n1536 = ~pi365 & ~n1534;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = pi362 & pi410;
  assign n1539 = ~n1537 & n1538;
  assign n1540 = ~pi362 & pi410;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = pi363 & n1541;
  assign n1543 = ~pi363 & ~n1541;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = pi322 & ~n1544;
  assign n1546 = ~n1531 & n1545;
  assign n1547 = ~pi322 & ~n1544;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = pi323 & n1548;
  assign n1550 = ~pi323 & ~n1548;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = pi282 & ~n1551;
  assign n1553 = ~n1525 & n1552;
  assign n1554 = ~pi282 & ~n1551;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = pi283 & n1555;
  assign n1557 = ~pi283 & ~n1555;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = pi242 & ~n1558;
  assign n1560 = ~n1519 & n1559;
  assign n1561 = ~pi242 & ~n1558;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = pi243 & n1562;
  assign n1564 = ~pi243 & ~n1562;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = pi202 & ~n1565;
  assign n1567 = ~n1513 & n1566;
  assign n1568 = ~pi202 & ~n1565;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = pi203 & n1569;
  assign n1571 = ~pi203 & ~n1569;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = pi162 & ~n1572;
  assign n1574 = ~n1507 & n1573;
  assign n1575 = ~pi162 & ~n1572;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = pi163 & n1576;
  assign n1578 = ~pi163 & ~n1576;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = pi122 & ~n1579;
  assign n1581 = ~n1501 & n1580;
  assign n1582 = ~pi122 & ~n1579;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = pi123 & n1583;
  assign n1585 = ~pi123 & ~n1583;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = pi082 & ~n1586;
  assign n1588 = ~n1495 & n1587;
  assign n1589 = ~pi082 & ~n1586;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = pi083 & n1590;
  assign n1592 = ~pi083 & ~n1590;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = pi042 & ~n1593;
  assign n1595 = ~n1489 & n1594;
  assign n1596 = ~pi042 & ~n1593;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = pi043 & n1597;
  assign n1599 = ~pi043 & ~n1597;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = pi000 & ~n1483;
  assign n1602 = ~n1600 & n1601;
  assign n1603 = ~pi000 & ~n1483;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = pi001 & n1604;
  assign n1606 = ~pi001 & ~n1604;
  assign po0 = n1605 | n1606;
endmodule


