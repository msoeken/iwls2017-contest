// Benchmark "trans_arith" written by ABC on Wed Apr 26 18:23:08 2017

module trans_arith ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825;
  assign n83 = pi40 & pi64;
  assign n84 = pi48 & ~pi64;
  assign n85 = ~n83 & ~n84;
  assign n86 = pi16 & pi24;
  assign n87 = n85 & n86;
  assign n88 = ~n85 & ~n86;
  assign n89 = ~n87 & ~n88;
  assign n90 = pi08 & pi64;
  assign n91 = pi32 & ~pi64;
  assign n92 = ~n90 & ~n91;
  assign n93 = pi00 & pi56;
  assign n94 = ~n92 & n93;
  assign n95 = n92 & ~n93;
  assign n96 = ~n94 & ~n95;
  assign po00 = ~n89 & n96;
  assign n98 = pi41 & pi64;
  assign n99 = pi49 & ~pi64;
  assign n100 = ~n98 & ~n99;
  assign n101 = pi17 & pi24;
  assign n102 = pi16 & pi25;
  assign n103 = n101 & n102;
  assign n104 = ~n101 & ~n102;
  assign n105 = ~n103 & ~n104;
  assign n106 = ~n100 & ~n105;
  assign n107 = n100 & n105;
  assign n108 = ~n106 & ~n107;
  assign n109 = ~n87 & n108;
  assign n110 = n87 & ~n108;
  assign n111 = ~n109 & ~n110;
  assign n112 = n96 & n111;
  assign n113 = pi09 & pi64;
  assign n114 = pi33 & ~pi64;
  assign n115 = ~n113 & ~n114;
  assign n116 = pi01 & pi56;
  assign n117 = pi00 & pi57;
  assign n118 = n116 & n117;
  assign n119 = ~n116 & ~n117;
  assign n120 = ~n118 & ~n119;
  assign n121 = ~n115 & n120;
  assign n122 = n115 & ~n120;
  assign n123 = ~n121 & ~n122;
  assign n124 = n94 & n123;
  assign n125 = ~n94 & ~n123;
  assign n126 = ~n124 & ~n125;
  assign n127 = ~n89 & n126;
  assign n128 = n112 & n127;
  assign n129 = ~n112 & ~n127;
  assign po01 = ~n128 & ~n129;
  assign n131 = ~n106 & ~n109;
  assign n132 = pi42 & pi64;
  assign n133 = pi50 & ~pi64;
  assign n134 = ~n132 & ~n133;
  assign n135 = pi18 & pi24;
  assign n136 = pi17 & pi25;
  assign n137 = n135 & n136;
  assign n138 = ~n135 & ~n136;
  assign n139 = ~n137 & ~n138;
  assign n140 = pi16 & pi26;
  assign n141 = n139 & n140;
  assign n142 = ~n139 & ~n140;
  assign n143 = ~n141 & ~n142;
  assign n144 = n103 & n143;
  assign n145 = ~n103 & ~n143;
  assign n146 = ~n144 & ~n145;
  assign n147 = ~n134 & ~n146;
  assign n148 = n134 & n146;
  assign n149 = ~n147 & ~n148;
  assign n150 = ~n131 & n149;
  assign n151 = n131 & ~n149;
  assign n152 = ~n150 & ~n151;
  assign n153 = n96 & n152;
  assign n154 = n111 & n126;
  assign n155 = n153 & n154;
  assign n156 = ~n153 & ~n154;
  assign n157 = ~n155 & ~n156;
  assign n158 = ~n121 & ~n124;
  assign n159 = pi10 & pi64;
  assign n160 = pi34 & ~pi64;
  assign n161 = ~n159 & ~n160;
  assign n162 = pi02 & pi56;
  assign n163 = pi01 & pi57;
  assign n164 = n162 & n163;
  assign n165 = ~n162 & ~n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = pi00 & pi58;
  assign n168 = n166 & n167;
  assign n169 = ~n166 & ~n167;
  assign n170 = ~n168 & ~n169;
  assign n171 = n118 & n170;
  assign n172 = ~n118 & ~n170;
  assign n173 = ~n171 & ~n172;
  assign n174 = ~n161 & n173;
  assign n175 = n161 & ~n173;
  assign n176 = ~n174 & ~n175;
  assign n177 = ~n158 & n176;
  assign n178 = n158 & ~n176;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n89 & n179;
  assign n181 = n157 & n180;
  assign n182 = ~n157 & ~n180;
  assign n183 = ~n181 & ~n182;
  assign n184 = n128 & n183;
  assign n185 = ~n128 & ~n183;
  assign po02 = ~n184 & ~n185;
  assign n187 = ~n181 & ~n184;
  assign n188 = ~n147 & ~n150;
  assign n189 = pi43 & pi64;
  assign n190 = pi51 & ~pi64;
  assign n191 = ~n189 & ~n190;
  assign n192 = ~n141 & ~n144;
  assign n193 = pi19 & pi24;
  assign n194 = pi18 & pi25;
  assign n195 = n193 & n194;
  assign n196 = ~n193 & ~n194;
  assign n197 = ~n195 & ~n196;
  assign n198 = pi17 & pi26;
  assign n199 = n197 & n198;
  assign n200 = ~n197 & ~n198;
  assign n201 = ~n199 & ~n200;
  assign n202 = n137 & n201;
  assign n203 = ~n137 & ~n201;
  assign n204 = ~n202 & ~n203;
  assign n205 = pi16 & pi27;
  assign n206 = n204 & n205;
  assign n207 = ~n204 & ~n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n192 & n208;
  assign n210 = n192 & ~n208;
  assign n211 = ~n209 & ~n210;
  assign n212 = ~n191 & ~n211;
  assign n213 = n191 & n211;
  assign n214 = ~n212 & ~n213;
  assign n215 = ~n188 & n214;
  assign n216 = n188 & ~n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = n96 & n217;
  assign n219 = n126 & n152;
  assign n220 = n218 & n219;
  assign n221 = ~n218 & ~n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = n111 & n179;
  assign n224 = n222 & n223;
  assign n225 = ~n222 & ~n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = n155 & n226;
  assign n228 = ~n155 & ~n226;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~n174 & ~n177;
  assign n231 = pi11 & pi64;
  assign n232 = pi35 & ~pi64;
  assign n233 = ~n231 & ~n232;
  assign n234 = ~n168 & ~n171;
  assign n235 = pi03 & pi56;
  assign n236 = pi02 & pi57;
  assign n237 = n235 & n236;
  assign n238 = ~n235 & ~n236;
  assign n239 = ~n237 & ~n238;
  assign n240 = pi01 & pi58;
  assign n241 = n239 & n240;
  assign n242 = ~n239 & ~n240;
  assign n243 = ~n241 & ~n242;
  assign n244 = n164 & n243;
  assign n245 = ~n164 & ~n243;
  assign n246 = ~n244 & ~n245;
  assign n247 = pi00 & pi59;
  assign n248 = n246 & n247;
  assign n249 = ~n246 & ~n247;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n234 & n250;
  assign n252 = n234 & ~n250;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~n233 & n253;
  assign n255 = n233 & ~n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = ~n230 & n256;
  assign n258 = n230 & ~n256;
  assign n259 = ~n257 & ~n258;
  assign n260 = ~n89 & n259;
  assign n261 = n229 & n260;
  assign n262 = ~n229 & ~n260;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n187 & n263;
  assign n265 = n187 & ~n263;
  assign po03 = ~n264 & ~n265;
  assign n267 = ~n261 & ~n264;
  assign n268 = ~n224 & ~n227;
  assign n269 = ~n212 & ~n215;
  assign n270 = pi44 & pi64;
  assign n271 = pi52 & ~pi64;
  assign n272 = ~n270 & ~n271;
  assign n273 = ~n206 & ~n209;
  assign n274 = ~n199 & ~n202;
  assign n275 = pi20 & pi24;
  assign n276 = pi19 & pi25;
  assign n277 = n275 & n276;
  assign n278 = ~n275 & ~n276;
  assign n279 = ~n277 & ~n278;
  assign n280 = pi18 & pi26;
  assign n281 = n279 & n280;
  assign n282 = ~n279 & ~n280;
  assign n283 = ~n281 & ~n282;
  assign n284 = n195 & n283;
  assign n285 = ~n195 & ~n283;
  assign n286 = ~n284 & ~n285;
  assign n287 = pi17 & pi27;
  assign n288 = n286 & n287;
  assign n289 = ~n286 & ~n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n274 & n290;
  assign n292 = n274 & ~n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = pi16 & pi28;
  assign n295 = n293 & n294;
  assign n296 = ~n293 & ~n294;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n273 & n297;
  assign n299 = n273 & ~n297;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~n272 & ~n300;
  assign n302 = n272 & n300;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n269 & n303;
  assign n305 = n269 & ~n303;
  assign n306 = ~n304 & ~n305;
  assign n307 = n96 & n306;
  assign n308 = n126 & n217;
  assign n309 = n307 & n308;
  assign n310 = ~n307 & ~n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = n152 & n179;
  assign n313 = n311 & n312;
  assign n314 = ~n311 & ~n312;
  assign n315 = ~n313 & ~n314;
  assign n316 = n220 & n315;
  assign n317 = ~n220 & ~n315;
  assign n318 = ~n316 & ~n317;
  assign n319 = n111 & n259;
  assign n320 = n318 & n319;
  assign n321 = ~n318 & ~n319;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~n268 & n322;
  assign n324 = n268 & ~n322;
  assign n325 = ~n323 & ~n324;
  assign n326 = ~n254 & ~n257;
  assign n327 = pi12 & pi64;
  assign n328 = pi36 & ~pi64;
  assign n329 = ~n327 & ~n328;
  assign n330 = ~n248 & ~n251;
  assign n331 = ~n241 & ~n244;
  assign n332 = pi04 & pi56;
  assign n333 = pi03 & pi57;
  assign n334 = n332 & n333;
  assign n335 = ~n332 & ~n333;
  assign n336 = ~n334 & ~n335;
  assign n337 = pi02 & pi58;
  assign n338 = n336 & n337;
  assign n339 = ~n336 & ~n337;
  assign n340 = ~n338 & ~n339;
  assign n341 = n237 & n340;
  assign n342 = ~n237 & ~n340;
  assign n343 = ~n341 & ~n342;
  assign n344 = pi01 & pi59;
  assign n345 = n343 & n344;
  assign n346 = ~n343 & ~n344;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~n331 & n347;
  assign n349 = n331 & ~n347;
  assign n350 = ~n348 & ~n349;
  assign n351 = pi00 & pi60;
  assign n352 = n350 & n351;
  assign n353 = ~n350 & ~n351;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~n330 & n354;
  assign n356 = n330 & ~n354;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n329 & n357;
  assign n359 = n329 & ~n357;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n326 & n360;
  assign n362 = n326 & ~n360;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~n89 & n363;
  assign n365 = n325 & n364;
  assign n366 = ~n325 & ~n364;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~n267 & n367;
  assign n369 = n267 & ~n367;
  assign po04 = ~n368 & ~n369;
  assign n371 = ~n365 & ~n368;
  assign n372 = ~n320 & ~n323;
  assign n373 = ~n313 & ~n316;
  assign n374 = ~n301 & ~n304;
  assign n375 = pi45 & pi64;
  assign n376 = pi53 & ~pi64;
  assign n377 = ~n375 & ~n376;
  assign n378 = ~n295 & ~n298;
  assign n379 = ~n288 & ~n291;
  assign n380 = ~n281 & ~n284;
  assign n381 = pi21 & pi24;
  assign n382 = pi20 & pi25;
  assign n383 = n381 & n382;
  assign n384 = ~n381 & ~n382;
  assign n385 = ~n383 & ~n384;
  assign n386 = pi19 & pi26;
  assign n387 = n385 & n386;
  assign n388 = ~n385 & ~n386;
  assign n389 = ~n387 & ~n388;
  assign n390 = n277 & n389;
  assign n391 = ~n277 & ~n389;
  assign n392 = ~n390 & ~n391;
  assign n393 = pi18 & pi27;
  assign n394 = n392 & n393;
  assign n395 = ~n392 & ~n393;
  assign n396 = ~n394 & ~n395;
  assign n397 = ~n380 & n396;
  assign n398 = n380 & ~n396;
  assign n399 = ~n397 & ~n398;
  assign n400 = pi17 & pi28;
  assign n401 = n399 & n400;
  assign n402 = ~n399 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n379 & n403;
  assign n405 = n379 & ~n403;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi16 & pi29;
  assign n408 = n406 & n407;
  assign n409 = ~n406 & ~n407;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~n378 & n410;
  assign n412 = n378 & ~n410;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~n377 & ~n413;
  assign n415 = n377 & n413;
  assign n416 = ~n414 & ~n415;
  assign n417 = ~n374 & n416;
  assign n418 = n374 & ~n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = n96 & n419;
  assign n421 = n126 & n306;
  assign n422 = n420 & n421;
  assign n423 = ~n420 & ~n421;
  assign n424 = ~n422 & ~n423;
  assign n425 = n179 & n217;
  assign n426 = n424 & n425;
  assign n427 = ~n424 & ~n425;
  assign n428 = ~n426 & ~n427;
  assign n429 = n309 & n428;
  assign n430 = ~n309 & ~n428;
  assign n431 = ~n429 & ~n430;
  assign n432 = n152 & n259;
  assign n433 = n431 & n432;
  assign n434 = ~n431 & ~n432;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~n373 & n435;
  assign n437 = n373 & ~n435;
  assign n438 = ~n436 & ~n437;
  assign n439 = n111 & n363;
  assign n440 = n438 & n439;
  assign n441 = ~n438 & ~n439;
  assign n442 = ~n440 & ~n441;
  assign n443 = ~n372 & n442;
  assign n444 = n372 & ~n442;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~n358 & ~n361;
  assign n447 = pi13 & pi64;
  assign n448 = pi37 & ~pi64;
  assign n449 = ~n447 & ~n448;
  assign n450 = ~n352 & ~n355;
  assign n451 = ~n345 & ~n348;
  assign n452 = ~n338 & ~n341;
  assign n453 = pi05 & pi56;
  assign n454 = pi04 & pi57;
  assign n455 = n453 & n454;
  assign n456 = ~n453 & ~n454;
  assign n457 = ~n455 & ~n456;
  assign n458 = pi03 & pi58;
  assign n459 = n457 & n458;
  assign n460 = ~n457 & ~n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = n334 & n461;
  assign n463 = ~n334 & ~n461;
  assign n464 = ~n462 & ~n463;
  assign n465 = pi02 & pi59;
  assign n466 = n464 & n465;
  assign n467 = ~n464 & ~n465;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~n452 & n468;
  assign n470 = n452 & ~n468;
  assign n471 = ~n469 & ~n470;
  assign n472 = pi01 & pi60;
  assign n473 = n471 & n472;
  assign n474 = ~n471 & ~n472;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n451 & n475;
  assign n477 = n451 & ~n475;
  assign n478 = ~n476 & ~n477;
  assign n479 = pi00 & pi61;
  assign n480 = n478 & n479;
  assign n481 = ~n478 & ~n479;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n450 & n482;
  assign n484 = n450 & ~n482;
  assign n485 = ~n483 & ~n484;
  assign n486 = ~n449 & n485;
  assign n487 = n449 & ~n485;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~n446 & n488;
  assign n490 = n446 & ~n488;
  assign n491 = ~n489 & ~n490;
  assign n492 = ~n89 & n491;
  assign n493 = n445 & n492;
  assign n494 = ~n445 & ~n492;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n371 & n495;
  assign n497 = n371 & ~n495;
  assign po05 = ~n496 & ~n497;
  assign n499 = ~n493 & ~n496;
  assign n500 = ~n440 & ~n443;
  assign n501 = ~n433 & ~n436;
  assign n502 = ~n426 & ~n429;
  assign n503 = ~n414 & ~n417;
  assign n504 = pi46 & pi64;
  assign n505 = pi54 & ~pi64;
  assign n506 = ~n504 & ~n505;
  assign n507 = ~n408 & ~n411;
  assign n508 = ~n401 & ~n404;
  assign n509 = ~n394 & ~n397;
  assign n510 = ~n387 & ~n390;
  assign n511 = pi22 & pi24;
  assign n512 = pi21 & pi25;
  assign n513 = n511 & n512;
  assign n514 = ~n511 & ~n512;
  assign n515 = ~n513 & ~n514;
  assign n516 = pi20 & pi26;
  assign n517 = n515 & n516;
  assign n518 = ~n515 & ~n516;
  assign n519 = ~n517 & ~n518;
  assign n520 = n383 & n519;
  assign n521 = ~n383 & ~n519;
  assign n522 = ~n520 & ~n521;
  assign n523 = pi19 & pi27;
  assign n524 = n522 & n523;
  assign n525 = ~n522 & ~n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~n510 & n526;
  assign n528 = n510 & ~n526;
  assign n529 = ~n527 & ~n528;
  assign n530 = pi18 & pi28;
  assign n531 = n529 & n530;
  assign n532 = ~n529 & ~n530;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~n509 & n533;
  assign n535 = n509 & ~n533;
  assign n536 = ~n534 & ~n535;
  assign n537 = pi17 & pi29;
  assign n538 = n536 & n537;
  assign n539 = ~n536 & ~n537;
  assign n540 = ~n538 & ~n539;
  assign n541 = ~n508 & n540;
  assign n542 = n508 & ~n540;
  assign n543 = ~n541 & ~n542;
  assign n544 = pi16 & pi30;
  assign n545 = n543 & n544;
  assign n546 = ~n543 & ~n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n507 & n547;
  assign n549 = n507 & ~n547;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~n506 & ~n550;
  assign n552 = n506 & n550;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n503 & n553;
  assign n555 = n503 & ~n553;
  assign n556 = ~n554 & ~n555;
  assign n557 = n96 & n556;
  assign n558 = n126 & n419;
  assign n559 = n557 & n558;
  assign n560 = ~n557 & ~n558;
  assign n561 = ~n559 & ~n560;
  assign n562 = n179 & n306;
  assign n563 = n561 & n562;
  assign n564 = ~n561 & ~n562;
  assign n565 = ~n563 & ~n564;
  assign n566 = n422 & n565;
  assign n567 = ~n422 & ~n565;
  assign n568 = ~n566 & ~n567;
  assign n569 = n217 & n259;
  assign n570 = n568 & n569;
  assign n571 = ~n568 & ~n569;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~n502 & n572;
  assign n574 = n502 & ~n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = n152 & n363;
  assign n577 = n575 & n576;
  assign n578 = ~n575 & ~n576;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n501 & n579;
  assign n581 = n501 & ~n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = n111 & n491;
  assign n584 = n582 & n583;
  assign n585 = ~n582 & ~n583;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n500 & n586;
  assign n588 = n500 & ~n586;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n486 & ~n489;
  assign n591 = pi14 & pi64;
  assign n592 = pi38 & ~pi64;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n480 & ~n483;
  assign n595 = ~n473 & ~n476;
  assign n596 = ~n466 & ~n469;
  assign n597 = ~n459 & ~n462;
  assign n598 = pi06 & pi56;
  assign n599 = pi05 & pi57;
  assign n600 = n598 & n599;
  assign n601 = ~n598 & ~n599;
  assign n602 = ~n600 & ~n601;
  assign n603 = pi04 & pi58;
  assign n604 = n602 & n603;
  assign n605 = ~n602 & ~n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = n455 & n606;
  assign n608 = ~n455 & ~n606;
  assign n609 = ~n607 & ~n608;
  assign n610 = pi03 & pi59;
  assign n611 = n609 & n610;
  assign n612 = ~n609 & ~n610;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n597 & n613;
  assign n615 = n597 & ~n613;
  assign n616 = ~n614 & ~n615;
  assign n617 = pi02 & pi60;
  assign n618 = n616 & n617;
  assign n619 = ~n616 & ~n617;
  assign n620 = ~n618 & ~n619;
  assign n621 = ~n596 & n620;
  assign n622 = n596 & ~n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = pi01 & pi61;
  assign n625 = n623 & n624;
  assign n626 = ~n623 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~n595 & n627;
  assign n629 = n595 & ~n627;
  assign n630 = ~n628 & ~n629;
  assign n631 = pi00 & pi62;
  assign n632 = n630 & n631;
  assign n633 = ~n630 & ~n631;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n594 & n634;
  assign n636 = n594 & ~n634;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~n593 & n637;
  assign n639 = n593 & ~n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n590 & n640;
  assign n642 = n590 & ~n640;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n89 & n643;
  assign n645 = n589 & n644;
  assign n646 = ~n589 & ~n644;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n499 & n647;
  assign n649 = n499 & ~n647;
  assign po06 = ~n648 & ~n649;
  assign n651 = ~n645 & ~n648;
  assign n652 = ~n584 & ~n587;
  assign n653 = ~n577 & ~n580;
  assign n654 = ~n570 & ~n573;
  assign n655 = ~n563 & ~n566;
  assign n656 = ~n551 & ~n554;
  assign n657 = pi47 & pi64;
  assign n658 = pi55 & ~pi64;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~n545 & ~n548;
  assign n661 = ~n538 & ~n541;
  assign n662 = ~n531 & ~n534;
  assign n663 = ~n524 & ~n527;
  assign n664 = ~n517 & ~n520;
  assign n665 = pi23 & pi24;
  assign n666 = pi22 & pi25;
  assign n667 = n665 & n666;
  assign n668 = ~n665 & ~n666;
  assign n669 = ~n667 & ~n668;
  assign n670 = pi21 & pi26;
  assign n671 = n669 & n670;
  assign n672 = ~n669 & ~n670;
  assign n673 = ~n671 & ~n672;
  assign n674 = n513 & n673;
  assign n675 = ~n513 & ~n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = pi20 & pi27;
  assign n678 = n676 & n677;
  assign n679 = ~n676 & ~n677;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~n664 & n680;
  assign n682 = n664 & ~n680;
  assign n683 = ~n681 & ~n682;
  assign n684 = pi19 & pi28;
  assign n685 = n683 & n684;
  assign n686 = ~n683 & ~n684;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n663 & n687;
  assign n689 = n663 & ~n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = pi18 & pi29;
  assign n692 = n690 & n691;
  assign n693 = ~n690 & ~n691;
  assign n694 = ~n692 & ~n693;
  assign n695 = ~n662 & n694;
  assign n696 = n662 & ~n694;
  assign n697 = ~n695 & ~n696;
  assign n698 = pi17 & pi30;
  assign n699 = n697 & n698;
  assign n700 = ~n697 & ~n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n661 & n701;
  assign n703 = n661 & ~n701;
  assign n704 = ~n702 & ~n703;
  assign n705 = pi16 & pi31;
  assign n706 = n704 & n705;
  assign n707 = ~n704 & ~n705;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n660 & n708;
  assign n710 = n660 & ~n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n659 & ~n711;
  assign n713 = n659 & n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n656 & n714;
  assign n716 = n656 & ~n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = n96 & n717;
  assign n719 = n126 & n556;
  assign n720 = n718 & n719;
  assign n721 = ~n718 & ~n719;
  assign n722 = ~n720 & ~n721;
  assign n723 = n179 & n419;
  assign n724 = n722 & n723;
  assign n725 = ~n722 & ~n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = n559 & n726;
  assign n728 = ~n559 & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = n259 & n306;
  assign n731 = n729 & n730;
  assign n732 = ~n729 & ~n730;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n655 & n733;
  assign n735 = n655 & ~n733;
  assign n736 = ~n734 & ~n735;
  assign n737 = n217 & n363;
  assign n738 = n736 & n737;
  assign n739 = ~n736 & ~n737;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n654 & n740;
  assign n742 = n654 & ~n740;
  assign n743 = ~n741 & ~n742;
  assign n744 = n152 & n491;
  assign n745 = n743 & n744;
  assign n746 = ~n743 & ~n744;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~n653 & n747;
  assign n749 = n653 & ~n747;
  assign n750 = ~n748 & ~n749;
  assign n751 = n111 & n643;
  assign n752 = n750 & n751;
  assign n753 = ~n750 & ~n751;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n652 & n754;
  assign n756 = n652 & ~n754;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n638 & ~n641;
  assign n759 = pi15 & pi64;
  assign n760 = pi39 & ~pi64;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~n632 & ~n635;
  assign n763 = ~n625 & ~n628;
  assign n764 = ~n618 & ~n621;
  assign n765 = ~n611 & ~n614;
  assign n766 = ~n604 & ~n607;
  assign n767 = pi07 & pi56;
  assign n768 = pi06 & pi57;
  assign n769 = n767 & n768;
  assign n770 = ~n767 & ~n768;
  assign n771 = ~n769 & ~n770;
  assign n772 = pi05 & pi58;
  assign n773 = n771 & n772;
  assign n774 = ~n771 & ~n772;
  assign n775 = ~n773 & ~n774;
  assign n776 = n600 & n775;
  assign n777 = ~n600 & ~n775;
  assign n778 = ~n776 & ~n777;
  assign n779 = pi04 & pi59;
  assign n780 = n778 & n779;
  assign n781 = ~n778 & ~n779;
  assign n782 = ~n780 & ~n781;
  assign n783 = ~n766 & n782;
  assign n784 = n766 & ~n782;
  assign n785 = ~n783 & ~n784;
  assign n786 = pi03 & pi60;
  assign n787 = n785 & n786;
  assign n788 = ~n785 & ~n786;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~n765 & n789;
  assign n791 = n765 & ~n789;
  assign n792 = ~n790 & ~n791;
  assign n793 = pi02 & pi61;
  assign n794 = n792 & n793;
  assign n795 = ~n792 & ~n793;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~n764 & n796;
  assign n798 = n764 & ~n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = pi01 & pi62;
  assign n801 = n799 & n800;
  assign n802 = ~n799 & ~n800;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n763 & n803;
  assign n805 = n763 & ~n803;
  assign n806 = ~n804 & ~n805;
  assign n807 = pi00 & pi63;
  assign n808 = n806 & n807;
  assign n809 = ~n806 & ~n807;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~n762 & n810;
  assign n812 = n762 & ~n810;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n761 & n813;
  assign n815 = n761 & ~n813;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~n758 & n816;
  assign n818 = n758 & ~n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n89 & n819;
  assign n821 = n757 & n820;
  assign n822 = ~n757 & ~n820;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~n651 & n823;
  assign n825 = n651 & ~n823;
  assign po07 = ~n824 & ~n825;
  assign po08 = 1'b0;
  assign po09 = 1'b0;
  assign po10 = 1'b0;
  assign po11 = 1'b0;
  assign po12 = 1'b0;
  assign po13 = 1'b0;
  assign po14 = 1'b0;
  assign po15 = 1'b0;
endmodule


