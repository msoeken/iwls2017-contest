// Benchmark "" written by ABC on Wed Apr 26 17:11:53 2017

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129;
  wire n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3090, n3091,
    n3093, n3094, n3096, n3097, n3099, n3100, n3102, n3103, n3105, n3106,
    n3108, n3109, n3111, n3112, n3114, n3115, n3117, n3118, n3120, n3121,
    n3123, n3124, n3126, n3127, n3129, n3130, n3132, n3133, n3135, n3136,
    n3138, n3139, n3141, n3142, n3144, n3145, n3147, n3148, n3150, n3151,
    n3153, n3154, n3156, n3157, n3159, n3160, n3162, n3163, n3165, n3166,
    n3168, n3169, n3171, n3172, n3174, n3175, n3177, n3178, n3180, n3181,
    n3183, n3184, n3186, n3187, n3189, n3190, n3192, n3193, n3195, n3196,
    n3198, n3199, n3201, n3202, n3204, n3205, n3207, n3208, n3210, n3211,
    n3213, n3214, n3216, n3217, n3219, n3220, n3222, n3223, n3225, n3226,
    n3228, n3229, n3231, n3232, n3234, n3235, n3237, n3238, n3240, n3241,
    n3243, n3244, n3246, n3247, n3249, n3250, n3252, n3253, n3255, n3256,
    n3258, n3259, n3261, n3262, n3264, n3265, n3267, n3268, n3270, n3271,
    n3273, n3274, n3276, n3277, n3279, n3280, n3282, n3283, n3285, n3286,
    n3288, n3289, n3291, n3292, n3294, n3295, n3297, n3298, n3300, n3301,
    n3303, n3304, n3306, n3307, n3309, n3310, n3312, n3313, n3315, n3316,
    n3318, n3319, n3321, n3322, n3324, n3325, n3327, n3328, n3330, n3331,
    n3333, n3334, n3336, n3337, n3339, n3340, n3342, n3343, n3345, n3346,
    n3348, n3349, n3351, n3352, n3354, n3355, n3357, n3358, n3360, n3361,
    n3363, n3364, n3366, n3367, n3369, n3370, n3372, n3373, n3375, n3376,
    n3378, n3379, n3381, n3382, n3384, n3385, n3387, n3388, n3390, n3391,
    n3393, n3394, n3396, n3397, n3399, n3400, n3402, n3403, n3405, n3406,
    n3408, n3409, n3411, n3412, n3414, n3415, n3417, n3418, n3420, n3421,
    n3423, n3424, n3426, n3427, n3429, n3430, n3432, n3433, n3435, n3436,
    n3438, n3439, n3441, n3442, n3444, n3445, n3447, n3448, n3450, n3451,
    n3453, n3454, n3456, n3457, n3459, n3460, n3462, n3463, n3465, n3466,
    n3468, n3469, n3472, n3473;
  assign n643 = ~pi383 & pi511;
  assign n644 = pi383 & ~pi511;
  assign n645 = ~pi381 & pi509;
  assign n646 = ~pi382 & pi510;
  assign n647 = ~n645 & ~n646;
  assign n648 = pi380 & ~pi508;
  assign n649 = pi381 & ~pi509;
  assign n650 = ~n648 & ~n649;
  assign n651 = n647 & ~n650;
  assign n652 = pi382 & ~pi510;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n644 & ~n653;
  assign n655 = pi379 & ~pi507;
  assign n656 = ~pi378 & pi506;
  assign n657 = ~pi379 & pi507;
  assign n658 = ~n656 & ~n657;
  assign n659 = pi378 & ~pi506;
  assign n660 = pi377 & ~pi505;
  assign n661 = ~pi377 & pi505;
  assign n662 = pi376 & ~pi504;
  assign n663 = ~n661 & n662;
  assign n664 = ~n659 & ~n660;
  assign n665 = ~n663 & n664;
  assign n666 = n658 & ~n665;
  assign n667 = pi375 & ~pi503;
  assign n668 = ~pi374 & pi502;
  assign n669 = ~pi375 & pi503;
  assign n670 = ~n668 & ~n669;
  assign n671 = pi374 & ~pi502;
  assign n672 = pi373 & ~pi501;
  assign n673 = ~pi373 & pi501;
  assign n674 = pi372 & ~pi500;
  assign n675 = ~n673 & n674;
  assign n676 = ~n671 & ~n672;
  assign n677 = ~n675 & n676;
  assign n678 = n670 & ~n677;
  assign n679 = pi371 & ~pi499;
  assign n680 = ~pi370 & pi498;
  assign n681 = ~pi371 & pi499;
  assign n682 = ~n680 & ~n681;
  assign n683 = pi370 & ~pi498;
  assign n684 = pi369 & ~pi497;
  assign n685 = ~pi369 & pi497;
  assign n686 = pi368 & ~pi496;
  assign n687 = ~n685 & n686;
  assign n688 = ~n683 & ~n684;
  assign n689 = ~n687 & n688;
  assign n690 = n682 & ~n689;
  assign n691 = pi367 & ~pi495;
  assign n692 = ~pi367 & pi495;
  assign n693 = ~pi366 & pi494;
  assign n694 = ~n692 & ~n693;
  assign n695 = pi366 & ~pi494;
  assign n696 = pi365 & ~pi493;
  assign n697 = ~pi365 & pi493;
  assign n698 = pi364 & ~pi492;
  assign n699 = ~n697 & n698;
  assign n700 = ~n695 & ~n696;
  assign n701 = ~n699 & n700;
  assign n702 = n694 & ~n701;
  assign n703 = pi363 & ~pi491;
  assign n704 = ~pi362 & pi490;
  assign n705 = ~pi363 & pi491;
  assign n706 = ~n704 & ~n705;
  assign n707 = pi362 & ~pi490;
  assign n708 = pi361 & ~pi489;
  assign n709 = ~pi361 & pi489;
  assign n710 = pi360 & ~pi488;
  assign n711 = ~n709 & n710;
  assign n712 = ~n707 & ~n708;
  assign n713 = ~n711 & n712;
  assign n714 = n706 & ~n713;
  assign n715 = pi359 & ~pi487;
  assign n716 = ~pi358 & pi486;
  assign n717 = ~pi359 & pi487;
  assign n718 = ~n716 & ~n717;
  assign n719 = pi358 & ~pi486;
  assign n720 = pi357 & ~pi485;
  assign n721 = ~pi357 & pi485;
  assign n722 = pi356 & ~pi484;
  assign n723 = ~n721 & n722;
  assign n724 = ~n719 & ~n720;
  assign n725 = ~n723 & n724;
  assign n726 = n718 & ~n725;
  assign n727 = pi355 & ~pi483;
  assign n728 = ~pi354 & pi482;
  assign n729 = ~pi355 & pi483;
  assign n730 = ~n728 & ~n729;
  assign n731 = pi354 & ~pi482;
  assign n732 = pi353 & ~pi481;
  assign n733 = ~pi353 & pi481;
  assign n734 = pi352 & ~pi480;
  assign n735 = ~n733 & n734;
  assign n736 = ~n731 & ~n732;
  assign n737 = ~n735 & n736;
  assign n738 = n730 & ~n737;
  assign n739 = pi351 & ~pi479;
  assign n740 = ~pi351 & pi479;
  assign n741 = ~pi350 & pi478;
  assign n742 = ~n740 & ~n741;
  assign n743 = pi350 & ~pi478;
  assign n744 = pi349 & ~pi477;
  assign n745 = ~pi349 & pi477;
  assign n746 = pi348 & ~pi476;
  assign n747 = ~n745 & n746;
  assign n748 = ~n743 & ~n744;
  assign n749 = ~n747 & n748;
  assign n750 = n742 & ~n749;
  assign n751 = ~pi346 & pi474;
  assign n752 = ~pi347 & pi475;
  assign n753 = ~n751 & ~n752;
  assign n754 = pi346 & ~pi474;
  assign n755 = pi345 & ~pi473;
  assign n756 = ~pi345 & pi473;
  assign n757 = pi344 & ~pi472;
  assign n758 = ~n756 & n757;
  assign n759 = ~n754 & ~n755;
  assign n760 = ~n758 & n759;
  assign n761 = n753 & ~n760;
  assign n762 = pi347 & ~pi475;
  assign n763 = pi343 & ~pi471;
  assign n764 = ~pi342 & pi470;
  assign n765 = ~pi343 & pi471;
  assign n766 = ~n764 & ~n765;
  assign n767 = pi342 & ~pi470;
  assign n768 = pi341 & ~pi469;
  assign n769 = ~pi341 & pi469;
  assign n770 = pi340 & ~pi468;
  assign n771 = ~n769 & n770;
  assign n772 = ~n767 & ~n768;
  assign n773 = ~n771 & n772;
  assign n774 = n766 & ~n773;
  assign n775 = pi339 & ~pi467;
  assign n776 = ~pi338 & pi466;
  assign n777 = ~pi339 & pi467;
  assign n778 = ~n776 & ~n777;
  assign n779 = pi338 & ~pi466;
  assign n780 = pi337 & ~pi465;
  assign n781 = ~pi337 & pi465;
  assign n782 = pi336 & ~pi464;
  assign n783 = ~n781 & n782;
  assign n784 = ~n779 & ~n780;
  assign n785 = ~n783 & n784;
  assign n786 = n778 & ~n785;
  assign n787 = pi335 & ~pi463;
  assign n788 = ~pi335 & pi463;
  assign n789 = ~pi334 & pi462;
  assign n790 = ~n788 & ~n789;
  assign n791 = pi334 & ~pi462;
  assign n792 = pi333 & ~pi461;
  assign n793 = ~pi333 & pi461;
  assign n794 = pi332 & ~pi460;
  assign n795 = ~n793 & n794;
  assign n796 = ~n791 & ~n792;
  assign n797 = ~n795 & n796;
  assign n798 = n790 & ~n797;
  assign n799 = ~pi330 & pi458;
  assign n800 = ~pi331 & pi459;
  assign n801 = ~n799 & ~n800;
  assign n802 = pi330 & ~pi458;
  assign n803 = pi329 & ~pi457;
  assign n804 = ~pi329 & pi457;
  assign n805 = pi328 & ~pi456;
  assign n806 = ~n804 & n805;
  assign n807 = ~n802 & ~n803;
  assign n808 = ~n806 & n807;
  assign n809 = n801 & ~n808;
  assign n810 = pi331 & ~pi459;
  assign n811 = pi323 & ~pi451;
  assign n812 = ~pi322 & pi450;
  assign n813 = ~pi314 & pi442;
  assign n814 = ~pi315 & pi443;
  assign n815 = ~n813 & ~n814;
  assign n816 = pi311 & ~pi439;
  assign n817 = ~pi310 & pi438;
  assign n818 = ~pi311 & pi439;
  assign n819 = ~n817 & ~n818;
  assign n820 = pi310 & ~pi438;
  assign n821 = ~pi309 & pi437;
  assign n822 = ~pi436 & ~n821;
  assign n823 = pi308 & n822;
  assign n824 = pi307 & ~pi435;
  assign n825 = ~pi306 & pi434;
  assign n826 = ~pi307 & pi435;
  assign n827 = ~n825 & ~n826;
  assign n828 = pi306 & ~pi434;
  assign n829 = pi305 & ~pi433;
  assign n830 = ~pi305 & pi433;
  assign n831 = pi304 & ~pi432;
  assign n832 = ~n830 & n831;
  assign n833 = ~n828 & ~n829;
  assign n834 = ~n832 & n833;
  assign n835 = n827 & ~n834;
  assign n836 = ~n824 & ~n835;
  assign n837 = pi308 & ~n821;
  assign n838 = ~n822 & ~n837;
  assign n839 = ~n836 & ~n838;
  assign n840 = pi309 & ~pi437;
  assign n841 = ~n820 & ~n840;
  assign n842 = ~n823 & n841;
  assign n843 = ~n839 & n842;
  assign n844 = n819 & ~n843;
  assign n845 = ~n816 & ~n844;
  assign n846 = n815 & ~n845;
  assign n847 = pi303 & ~pi431;
  assign n848 = ~pi302 & pi430;
  assign n849 = ~pi303 & pi431;
  assign n850 = ~n848 & ~n849;
  assign n851 = ~pi301 & pi429;
  assign n852 = ~pi428 & ~n851;
  assign n853 = pi300 & n852;
  assign n854 = pi299 & ~pi427;
  assign n855 = ~pi298 & pi426;
  assign n856 = ~pi299 & pi427;
  assign n857 = ~n855 & ~n856;
  assign n858 = pi298 & ~pi426;
  assign n859 = pi297 & ~pi425;
  assign n860 = ~pi297 & pi425;
  assign n861 = pi296 & ~pi424;
  assign n862 = ~n860 & n861;
  assign n863 = ~n858 & ~n859;
  assign n864 = ~n862 & n863;
  assign n865 = n857 & ~n864;
  assign n866 = ~n854 & ~n865;
  assign n867 = pi300 & ~n851;
  assign n868 = ~n852 & ~n867;
  assign n869 = ~n866 & ~n868;
  assign n870 = pi301 & ~pi429;
  assign n871 = pi302 & ~pi430;
  assign n872 = ~n870 & ~n871;
  assign n873 = ~n853 & n872;
  assign n874 = ~n869 & n873;
  assign n875 = n850 & ~n874;
  assign n876 = ~pi279 & pi407;
  assign n877 = ~pi280 & pi408;
  assign n878 = pi278 & ~pi406;
  assign n879 = pi279 & ~pi407;
  assign n880 = ~pi278 & pi406;
  assign n881 = pi277 & ~pi405;
  assign n882 = ~pi277 & pi405;
  assign n883 = pi276 & ~pi404;
  assign n884 = ~pi276 & pi404;
  assign n885 = pi275 & ~pi403;
  assign n886 = ~pi275 & pi403;
  assign n887 = pi274 & ~pi402;
  assign n888 = ~pi274 & pi402;
  assign n889 = pi273 & ~pi401;
  assign n890 = ~pi273 & pi401;
  assign n891 = pi272 & ~pi400;
  assign n892 = ~pi272 & pi400;
  assign n893 = pi271 & ~pi399;
  assign n894 = ~pi271 & pi399;
  assign n895 = pi270 & ~pi398;
  assign n896 = ~pi270 & pi398;
  assign n897 = pi269 & ~pi397;
  assign n898 = ~pi269 & pi397;
  assign n899 = pi268 & ~pi396;
  assign n900 = ~pi268 & pi396;
  assign n901 = pi267 & ~pi395;
  assign n902 = ~pi267 & pi395;
  assign n903 = pi266 & ~pi394;
  assign n904 = ~pi266 & pi394;
  assign n905 = pi265 & ~pi393;
  assign n906 = ~pi265 & pi393;
  assign n907 = pi264 & ~pi392;
  assign n908 = ~pi264 & pi392;
  assign n909 = pi263 & ~pi391;
  assign n910 = ~pi263 & pi391;
  assign n911 = pi262 & ~pi390;
  assign n912 = ~pi262 & pi390;
  assign n913 = pi261 & ~pi389;
  assign n914 = ~pi261 & pi389;
  assign n915 = pi260 & ~pi388;
  assign n916 = ~pi260 & pi388;
  assign n917 = pi259 & ~pi387;
  assign n918 = ~pi259 & pi387;
  assign n919 = pi258 & ~pi386;
  assign n920 = ~pi258 & pi386;
  assign n921 = pi257 & ~pi385;
  assign n922 = ~pi257 & pi385;
  assign n923 = pi256 & ~pi384;
  assign n924 = ~n922 & n923;
  assign n925 = ~n921 & ~n924;
  assign n926 = ~n920 & ~n925;
  assign n927 = ~n919 & ~n926;
  assign n928 = ~n918 & ~n927;
  assign n929 = ~n917 & ~n928;
  assign n930 = ~n916 & ~n929;
  assign n931 = ~n915 & ~n930;
  assign n932 = ~n914 & ~n931;
  assign n933 = ~n913 & ~n932;
  assign n934 = ~n912 & ~n933;
  assign n935 = ~n911 & ~n934;
  assign n936 = ~n910 & ~n935;
  assign n937 = ~n909 & ~n936;
  assign n938 = ~n908 & ~n937;
  assign n939 = ~n907 & ~n938;
  assign n940 = ~n906 & ~n939;
  assign n941 = ~n905 & ~n940;
  assign n942 = ~n904 & ~n941;
  assign n943 = ~n903 & ~n942;
  assign n944 = ~n902 & ~n943;
  assign n945 = ~n901 & ~n944;
  assign n946 = ~n900 & ~n945;
  assign n947 = ~n899 & ~n946;
  assign n948 = ~n898 & ~n947;
  assign n949 = ~n897 & ~n948;
  assign n950 = ~n896 & ~n949;
  assign n951 = ~n895 & ~n950;
  assign n952 = ~n894 & ~n951;
  assign n953 = ~n893 & ~n952;
  assign n954 = ~n892 & ~n953;
  assign n955 = ~n891 & ~n954;
  assign n956 = ~n890 & ~n955;
  assign n957 = ~n889 & ~n956;
  assign n958 = ~n888 & ~n957;
  assign n959 = ~n887 & ~n958;
  assign n960 = ~n886 & ~n959;
  assign n961 = ~n885 & ~n960;
  assign n962 = ~n884 & ~n961;
  assign n963 = ~n883 & ~n962;
  assign n964 = ~n882 & ~n963;
  assign n965 = ~n881 & ~n964;
  assign n966 = ~n880 & ~n965;
  assign n967 = ~n878 & ~n879;
  assign n968 = ~n966 & n967;
  assign n969 = ~n876 & ~n877;
  assign n970 = ~n968 & n969;
  assign n971 = pi280 & ~pi408;
  assign n972 = pi281 & ~pi409;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n970 & n973;
  assign n975 = ~pi281 & pi409;
  assign n976 = ~pi282 & pi410;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n974 & n977;
  assign n979 = pi282 & ~pi410;
  assign n980 = pi283 & ~pi411;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n978 & n981;
  assign n983 = ~pi283 & pi411;
  assign n984 = ~pi284 & pi412;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~n982 & n985;
  assign n987 = pi284 & ~pi412;
  assign n988 = pi285 & ~pi413;
  assign n989 = ~n987 & ~n988;
  assign n990 = ~n986 & n989;
  assign n991 = ~pi285 & pi413;
  assign n992 = ~pi286 & pi414;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n990 & n993;
  assign n995 = pi286 & ~pi414;
  assign n996 = pi287 & ~pi415;
  assign n997 = ~n995 & ~n996;
  assign n998 = ~n994 & n997;
  assign n999 = ~pi292 & pi420;
  assign n1000 = ~pi290 & pi418;
  assign n1001 = ~pi291 & pi419;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~pi287 & pi415;
  assign n1004 = ~pi288 & pi416;
  assign n1005 = ~pi289 & pi417;
  assign n1006 = ~pi293 & pi421;
  assign n1007 = ~pi295 & pi423;
  assign n1008 = ~pi294 & pi422;
  assign n1009 = ~n1006 & ~n1007;
  assign n1010 = ~n1008 & n1009;
  assign n1011 = ~n999 & ~n1003;
  assign n1012 = ~n1004 & ~n1005;
  assign n1013 = n1011 & n1012;
  assign n1014 = n1002 & n1013;
  assign n1015 = n1010 & n1014;
  assign n1016 = ~n998 & n1015;
  assign n1017 = pi294 & ~pi422;
  assign n1018 = ~n1007 & n1017;
  assign n1019 = pi295 & ~pi423;
  assign n1020 = pi293 & ~pi421;
  assign n1021 = pi292 & ~pi420;
  assign n1022 = pi291 & ~pi419;
  assign n1023 = pi290 & ~pi418;
  assign n1024 = pi289 & ~pi417;
  assign n1025 = pi288 & ~pi416;
  assign n1026 = ~n1005 & n1025;
  assign n1027 = ~n1023 & ~n1024;
  assign n1028 = ~n1026 & n1027;
  assign n1029 = n1002 & ~n1028;
  assign n1030 = ~n1022 & ~n1029;
  assign n1031 = ~n999 & ~n1030;
  assign n1032 = ~n1020 & ~n1021;
  assign n1033 = ~n1031 & n1032;
  assign n1034 = n1010 & ~n1033;
  assign n1035 = ~n1018 & ~n1019;
  assign n1036 = ~n1034 & n1035;
  assign n1037 = ~n1016 & n1036;
  assign n1038 = ~pi296 & pi424;
  assign n1039 = ~n860 & ~n1038;
  assign n1040 = n850 & n1039;
  assign n1041 = n857 & n1040;
  assign n1042 = ~n868 & n1041;
  assign n1043 = ~n1037 & n1042;
  assign n1044 = ~n847 & ~n875;
  assign n1045 = ~n1043 & n1044;
  assign n1046 = ~pi304 & pi432;
  assign n1047 = ~n830 & ~n1046;
  assign n1048 = n819 & n1047;
  assign n1049 = n827 & n1048;
  assign n1050 = ~n838 & n1049;
  assign n1051 = ~n1045 & n1050;
  assign n1052 = ~n846 & ~n1051;
  assign n1053 = ~pi312 & pi440;
  assign n1054 = ~pi316 & pi444;
  assign n1055 = ~pi313 & pi441;
  assign n1056 = ~pi317 & pi445;
  assign n1057 = ~pi319 & pi447;
  assign n1058 = ~pi318 & pi446;
  assign n1059 = ~n1056 & ~n1057;
  assign n1060 = ~n1058 & n1059;
  assign n1061 = ~n1053 & ~n1054;
  assign n1062 = ~n1055 & n1061;
  assign n1063 = n815 & n1062;
  assign n1064 = n1060 & n1063;
  assign n1065 = ~n1052 & n1064;
  assign n1066 = pi318 & ~pi446;
  assign n1067 = ~n1057 & n1066;
  assign n1068 = pi319 & ~pi447;
  assign n1069 = pi317 & ~pi445;
  assign n1070 = pi316 & ~pi444;
  assign n1071 = pi315 & ~pi443;
  assign n1072 = pi314 & ~pi442;
  assign n1073 = pi313 & ~pi441;
  assign n1074 = pi312 & ~pi440;
  assign n1075 = ~n1055 & n1074;
  assign n1076 = ~n1072 & ~n1073;
  assign n1077 = ~n1075 & n1076;
  assign n1078 = n815 & ~n1077;
  assign n1079 = ~n1071 & ~n1078;
  assign n1080 = ~n1054 & ~n1079;
  assign n1081 = ~n1069 & ~n1070;
  assign n1082 = ~n1080 & n1081;
  assign n1083 = n1060 & ~n1082;
  assign n1084 = ~n1067 & ~n1068;
  assign n1085 = ~n1083 & n1084;
  assign n1086 = ~n1065 & n1085;
  assign n1087 = ~pi321 & pi449;
  assign n1088 = ~pi320 & pi448;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n1086 & n1089;
  assign n1091 = pi322 & ~pi450;
  assign n1092 = pi321 & ~pi449;
  assign n1093 = pi320 & ~pi448;
  assign n1094 = ~n1087 & n1093;
  assign n1095 = ~n1091 & ~n1092;
  assign n1096 = ~n1094 & n1095;
  assign n1097 = ~n1090 & n1096;
  assign n1098 = ~n812 & ~n1097;
  assign n1099 = ~n811 & ~n1098;
  assign n1100 = ~pi325 & pi453;
  assign n1101 = ~pi324 & pi452;
  assign n1102 = ~pi326 & pi454;
  assign n1103 = ~pi327 & pi455;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~pi323 & pi451;
  assign n1106 = ~n1100 & ~n1101;
  assign n1107 = ~n1105 & n1106;
  assign n1108 = n1104 & n1107;
  assign n1109 = ~n1099 & n1108;
  assign n1110 = pi327 & ~pi455;
  assign n1111 = pi326 & ~pi454;
  assign n1112 = pi325 & ~pi453;
  assign n1113 = pi324 & ~pi452;
  assign n1114 = ~n1100 & n1113;
  assign n1115 = ~n1111 & ~n1112;
  assign n1116 = ~n1114 & n1115;
  assign n1117 = n1104 & ~n1116;
  assign n1118 = ~n1110 & ~n1117;
  assign n1119 = ~n1109 & n1118;
  assign n1120 = ~pi328 & pi456;
  assign n1121 = ~n804 & ~n1120;
  assign n1122 = n801 & n1121;
  assign n1123 = ~n1119 & n1122;
  assign n1124 = ~n809 & ~n810;
  assign n1125 = ~n1123 & n1124;
  assign n1126 = ~pi332 & pi460;
  assign n1127 = ~n793 & ~n1126;
  assign n1128 = n790 & n1127;
  assign n1129 = ~n1125 & n1128;
  assign n1130 = ~n787 & ~n798;
  assign n1131 = ~n1129 & n1130;
  assign n1132 = ~pi336 & pi464;
  assign n1133 = ~n781 & ~n1132;
  assign n1134 = n778 & n1133;
  assign n1135 = ~n1131 & n1134;
  assign n1136 = ~n775 & ~n786;
  assign n1137 = ~n1135 & n1136;
  assign n1138 = ~pi340 & pi468;
  assign n1139 = ~n769 & ~n1138;
  assign n1140 = n766 & n1139;
  assign n1141 = ~n1137 & n1140;
  assign n1142 = ~n763 & ~n774;
  assign n1143 = ~n1141 & n1142;
  assign n1144 = ~pi344 & pi472;
  assign n1145 = ~n756 & ~n1144;
  assign n1146 = n753 & n1145;
  assign n1147 = ~n1143 & n1146;
  assign n1148 = ~n761 & ~n762;
  assign n1149 = ~n1147 & n1148;
  assign n1150 = ~pi348 & pi476;
  assign n1151 = ~n745 & ~n1150;
  assign n1152 = n742 & n1151;
  assign n1153 = ~n1149 & n1152;
  assign n1154 = ~n739 & ~n750;
  assign n1155 = ~n1153 & n1154;
  assign n1156 = ~pi352 & pi480;
  assign n1157 = ~n733 & ~n1156;
  assign n1158 = n730 & n1157;
  assign n1159 = ~n1155 & n1158;
  assign n1160 = ~n727 & ~n738;
  assign n1161 = ~n1159 & n1160;
  assign n1162 = ~pi356 & pi484;
  assign n1163 = ~n721 & ~n1162;
  assign n1164 = n718 & n1163;
  assign n1165 = ~n1161 & n1164;
  assign n1166 = ~n715 & ~n726;
  assign n1167 = ~n1165 & n1166;
  assign n1168 = ~pi360 & pi488;
  assign n1169 = ~n709 & ~n1168;
  assign n1170 = n706 & n1169;
  assign n1171 = ~n1167 & n1170;
  assign n1172 = ~n703 & ~n714;
  assign n1173 = ~n1171 & n1172;
  assign n1174 = ~pi364 & pi492;
  assign n1175 = ~n697 & ~n1174;
  assign n1176 = n694 & n1175;
  assign n1177 = ~n1173 & n1176;
  assign n1178 = ~n691 & ~n702;
  assign n1179 = ~n1177 & n1178;
  assign n1180 = ~pi368 & pi496;
  assign n1181 = ~n685 & ~n1180;
  assign n1182 = n682 & n1181;
  assign n1183 = ~n1179 & n1182;
  assign n1184 = ~n679 & ~n690;
  assign n1185 = ~n1183 & n1184;
  assign n1186 = ~pi372 & pi500;
  assign n1187 = ~n673 & ~n1186;
  assign n1188 = n670 & n1187;
  assign n1189 = ~n1185 & n1188;
  assign n1190 = ~n667 & ~n678;
  assign n1191 = ~n1189 & n1190;
  assign n1192 = ~pi376 & pi504;
  assign n1193 = ~n661 & ~n1192;
  assign n1194 = n658 & n1193;
  assign n1195 = ~n1191 & n1194;
  assign n1196 = ~n655 & ~n666;
  assign n1197 = ~n1195 & n1196;
  assign n1198 = ~pi380 & pi508;
  assign n1199 = ~n644 & ~n1198;
  assign n1200 = n647 & n1199;
  assign n1201 = ~n1197 & n1200;
  assign n1202 = ~n643 & ~n654;
  assign n1203 = ~n1201 & n1202;
  assign n1204 = pi256 & ~n1203;
  assign n1205 = pi384 & n1203;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = pi127 & ~pi255;
  assign n1208 = ~pi125 & pi253;
  assign n1209 = ~pi126 & pi254;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = pi124 & ~pi252;
  assign n1212 = pi125 & ~pi253;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = n1210 & ~n1213;
  assign n1215 = pi126 & ~pi254;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1207 & ~n1216;
  assign n1218 = ~pi127 & pi255;
  assign n1219 = pi123 & ~pi251;
  assign n1220 = ~pi122 & pi250;
  assign n1221 = ~pi123 & pi251;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = pi122 & ~pi250;
  assign n1224 = pi121 & ~pi249;
  assign n1225 = ~pi121 & pi249;
  assign n1226 = pi120 & ~pi248;
  assign n1227 = ~n1225 & n1226;
  assign n1228 = ~n1223 & ~n1224;
  assign n1229 = ~n1227 & n1228;
  assign n1230 = n1222 & ~n1229;
  assign n1231 = pi119 & ~pi247;
  assign n1232 = ~pi118 & pi246;
  assign n1233 = ~pi119 & pi247;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = pi118 & ~pi246;
  assign n1236 = pi117 & ~pi245;
  assign n1237 = ~pi117 & pi245;
  assign n1238 = pi116 & ~pi244;
  assign n1239 = ~n1237 & n1238;
  assign n1240 = ~n1235 & ~n1236;
  assign n1241 = ~n1239 & n1240;
  assign n1242 = n1234 & ~n1241;
  assign n1243 = pi115 & ~pi243;
  assign n1244 = ~pi114 & pi242;
  assign n1245 = ~pi115 & pi243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = pi114 & ~pi242;
  assign n1248 = pi113 & ~pi241;
  assign n1249 = ~pi113 & pi241;
  assign n1250 = pi112 & ~pi240;
  assign n1251 = ~n1249 & n1250;
  assign n1252 = ~n1247 & ~n1248;
  assign n1253 = ~n1251 & n1252;
  assign n1254 = n1246 & ~n1253;
  assign n1255 = pi111 & ~pi239;
  assign n1256 = ~pi111 & pi239;
  assign n1257 = ~pi110 & pi238;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = pi110 & ~pi238;
  assign n1260 = pi109 & ~pi237;
  assign n1261 = ~pi109 & pi237;
  assign n1262 = pi108 & ~pi236;
  assign n1263 = ~n1261 & n1262;
  assign n1264 = ~n1259 & ~n1260;
  assign n1265 = ~n1263 & n1264;
  assign n1266 = n1258 & ~n1265;
  assign n1267 = pi107 & ~pi235;
  assign n1268 = ~pi106 & pi234;
  assign n1269 = ~pi107 & pi235;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = pi106 & ~pi234;
  assign n1272 = pi105 & ~pi233;
  assign n1273 = ~pi105 & pi233;
  assign n1274 = pi104 & ~pi232;
  assign n1275 = ~n1273 & n1274;
  assign n1276 = ~n1271 & ~n1272;
  assign n1277 = ~n1275 & n1276;
  assign n1278 = n1270 & ~n1277;
  assign n1279 = pi103 & ~pi231;
  assign n1280 = ~pi102 & pi230;
  assign n1281 = ~pi103 & pi231;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = pi102 & ~pi230;
  assign n1284 = pi101 & ~pi229;
  assign n1285 = ~pi101 & pi229;
  assign n1286 = pi100 & ~pi228;
  assign n1287 = ~n1285 & n1286;
  assign n1288 = ~n1283 & ~n1284;
  assign n1289 = ~n1287 & n1288;
  assign n1290 = n1282 & ~n1289;
  assign n1291 = pi099 & ~pi227;
  assign n1292 = ~pi098 & pi226;
  assign n1293 = ~pi099 & pi227;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = pi098 & ~pi226;
  assign n1296 = pi097 & ~pi225;
  assign n1297 = ~pi097 & pi225;
  assign n1298 = pi096 & ~pi224;
  assign n1299 = ~n1297 & n1298;
  assign n1300 = ~n1295 & ~n1296;
  assign n1301 = ~n1299 & n1300;
  assign n1302 = n1294 & ~n1301;
  assign n1303 = pi095 & ~pi223;
  assign n1304 = ~pi095 & pi223;
  assign n1305 = ~pi094 & pi222;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = pi094 & ~pi222;
  assign n1308 = pi093 & ~pi221;
  assign n1309 = ~pi093 & pi221;
  assign n1310 = pi092 & ~pi220;
  assign n1311 = ~n1309 & n1310;
  assign n1312 = ~n1307 & ~n1308;
  assign n1313 = ~n1311 & n1312;
  assign n1314 = n1306 & ~n1313;
  assign n1315 = ~pi090 & pi218;
  assign n1316 = ~pi091 & pi219;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = pi090 & ~pi218;
  assign n1319 = pi089 & ~pi217;
  assign n1320 = ~pi089 & pi217;
  assign n1321 = pi088 & ~pi216;
  assign n1322 = ~n1320 & n1321;
  assign n1323 = ~n1318 & ~n1319;
  assign n1324 = ~n1322 & n1323;
  assign n1325 = n1317 & ~n1324;
  assign n1326 = pi091 & ~pi219;
  assign n1327 = pi087 & ~pi215;
  assign n1328 = ~pi086 & pi214;
  assign n1329 = ~pi087 & pi215;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = pi086 & ~pi214;
  assign n1332 = pi085 & ~pi213;
  assign n1333 = ~pi085 & pi213;
  assign n1334 = pi084 & ~pi212;
  assign n1335 = ~n1333 & n1334;
  assign n1336 = ~n1331 & ~n1332;
  assign n1337 = ~n1335 & n1336;
  assign n1338 = n1330 & ~n1337;
  assign n1339 = pi083 & ~pi211;
  assign n1340 = ~pi082 & pi210;
  assign n1341 = ~pi083 & pi211;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = pi082 & ~pi210;
  assign n1344 = pi081 & ~pi209;
  assign n1345 = ~pi081 & pi209;
  assign n1346 = pi080 & ~pi208;
  assign n1347 = ~n1345 & n1346;
  assign n1348 = ~n1343 & ~n1344;
  assign n1349 = ~n1347 & n1348;
  assign n1350 = n1342 & ~n1349;
  assign n1351 = pi079 & ~pi207;
  assign n1352 = ~pi079 & pi207;
  assign n1353 = ~pi078 & pi206;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = pi078 & ~pi206;
  assign n1356 = pi077 & ~pi205;
  assign n1357 = ~pi077 & pi205;
  assign n1358 = pi076 & ~pi204;
  assign n1359 = ~n1357 & n1358;
  assign n1360 = ~n1355 & ~n1356;
  assign n1361 = ~n1359 & n1360;
  assign n1362 = n1354 & ~n1361;
  assign n1363 = ~pi074 & pi202;
  assign n1364 = ~pi075 & pi203;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = pi074 & ~pi202;
  assign n1367 = pi073 & ~pi201;
  assign n1368 = ~pi073 & pi201;
  assign n1369 = pi072 & ~pi200;
  assign n1370 = ~n1368 & n1369;
  assign n1371 = ~n1366 & ~n1367;
  assign n1372 = ~n1370 & n1371;
  assign n1373 = n1365 & ~n1372;
  assign n1374 = pi075 & ~pi203;
  assign n1375 = pi067 & ~pi195;
  assign n1376 = ~pi066 & pi194;
  assign n1377 = ~pi058 & pi186;
  assign n1378 = ~pi059 & pi187;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = pi055 & ~pi183;
  assign n1381 = ~pi054 & pi182;
  assign n1382 = ~pi055 & pi183;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = pi054 & ~pi182;
  assign n1385 = ~pi053 & pi181;
  assign n1386 = ~pi180 & ~n1385;
  assign n1387 = pi052 & n1386;
  assign n1388 = pi051 & ~pi179;
  assign n1389 = ~pi050 & pi178;
  assign n1390 = ~pi051 & pi179;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = pi050 & ~pi178;
  assign n1393 = pi049 & ~pi177;
  assign n1394 = ~pi049 & pi177;
  assign n1395 = pi048 & ~pi176;
  assign n1396 = ~n1394 & n1395;
  assign n1397 = ~n1392 & ~n1393;
  assign n1398 = ~n1396 & n1397;
  assign n1399 = n1391 & ~n1398;
  assign n1400 = ~n1388 & ~n1399;
  assign n1401 = pi052 & ~n1385;
  assign n1402 = ~n1386 & ~n1401;
  assign n1403 = ~n1400 & ~n1402;
  assign n1404 = pi053 & ~pi181;
  assign n1405 = ~n1384 & ~n1404;
  assign n1406 = ~n1387 & n1405;
  assign n1407 = ~n1403 & n1406;
  assign n1408 = n1383 & ~n1407;
  assign n1409 = ~n1380 & ~n1408;
  assign n1410 = n1379 & ~n1409;
  assign n1411 = pi047 & ~pi175;
  assign n1412 = ~pi046 & pi174;
  assign n1413 = ~pi047 & pi175;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~pi045 & pi173;
  assign n1416 = ~pi172 & ~n1415;
  assign n1417 = pi044 & n1416;
  assign n1418 = pi043 & ~pi171;
  assign n1419 = ~pi042 & pi170;
  assign n1420 = ~pi043 & pi171;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = pi042 & ~pi170;
  assign n1423 = pi041 & ~pi169;
  assign n1424 = ~pi041 & pi169;
  assign n1425 = pi040 & ~pi168;
  assign n1426 = ~n1424 & n1425;
  assign n1427 = ~n1422 & ~n1423;
  assign n1428 = ~n1426 & n1427;
  assign n1429 = n1421 & ~n1428;
  assign n1430 = ~n1418 & ~n1429;
  assign n1431 = pi044 & ~n1415;
  assign n1432 = ~n1416 & ~n1431;
  assign n1433 = ~n1430 & ~n1432;
  assign n1434 = pi045 & ~pi173;
  assign n1435 = pi046 & ~pi174;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n1417 & n1436;
  assign n1438 = ~n1433 & n1437;
  assign n1439 = n1414 & ~n1438;
  assign n1440 = ~pi023 & pi151;
  assign n1441 = ~pi024 & pi152;
  assign n1442 = pi022 & ~pi150;
  assign n1443 = pi023 & ~pi151;
  assign n1444 = ~pi022 & pi150;
  assign n1445 = pi021 & ~pi149;
  assign n1446 = ~pi021 & pi149;
  assign n1447 = pi020 & ~pi148;
  assign n1448 = ~pi020 & pi148;
  assign n1449 = pi019 & ~pi147;
  assign n1450 = ~pi019 & pi147;
  assign n1451 = pi018 & ~pi146;
  assign n1452 = ~pi018 & pi146;
  assign n1453 = pi017 & ~pi145;
  assign n1454 = ~pi017 & pi145;
  assign n1455 = pi016 & ~pi144;
  assign n1456 = ~pi016 & pi144;
  assign n1457 = pi015 & ~pi143;
  assign n1458 = ~pi015 & pi143;
  assign n1459 = pi014 & ~pi142;
  assign n1460 = ~pi014 & pi142;
  assign n1461 = pi013 & ~pi141;
  assign n1462 = ~pi013 & pi141;
  assign n1463 = pi012 & ~pi140;
  assign n1464 = ~pi012 & pi140;
  assign n1465 = pi011 & ~pi139;
  assign n1466 = ~pi011 & pi139;
  assign n1467 = pi010 & ~pi138;
  assign n1468 = ~pi010 & pi138;
  assign n1469 = pi009 & ~pi137;
  assign n1470 = ~pi009 & pi137;
  assign n1471 = pi008 & ~pi136;
  assign n1472 = ~pi008 & pi136;
  assign n1473 = pi007 & ~pi135;
  assign n1474 = ~pi007 & pi135;
  assign n1475 = pi006 & ~pi134;
  assign n1476 = ~pi006 & pi134;
  assign n1477 = pi005 & ~pi133;
  assign n1478 = ~pi005 & pi133;
  assign n1479 = pi004 & ~pi132;
  assign n1480 = ~pi004 & pi132;
  assign n1481 = pi003 & ~pi131;
  assign n1482 = ~pi003 & pi131;
  assign n1483 = pi002 & ~pi130;
  assign n1484 = ~pi002 & pi130;
  assign n1485 = pi001 & ~pi129;
  assign n1486 = ~pi001 & pi129;
  assign n1487 = pi000 & ~pi128;
  assign n1488 = ~n1486 & n1487;
  assign n1489 = ~n1485 & ~n1488;
  assign n1490 = ~n1484 & ~n1489;
  assign n1491 = ~n1483 & ~n1490;
  assign n1492 = ~n1482 & ~n1491;
  assign n1493 = ~n1481 & ~n1492;
  assign n1494 = ~n1480 & ~n1493;
  assign n1495 = ~n1479 & ~n1494;
  assign n1496 = ~n1478 & ~n1495;
  assign n1497 = ~n1477 & ~n1496;
  assign n1498 = ~n1476 & ~n1497;
  assign n1499 = ~n1475 & ~n1498;
  assign n1500 = ~n1474 & ~n1499;
  assign n1501 = ~n1473 & ~n1500;
  assign n1502 = ~n1472 & ~n1501;
  assign n1503 = ~n1471 & ~n1502;
  assign n1504 = ~n1470 & ~n1503;
  assign n1505 = ~n1469 & ~n1504;
  assign n1506 = ~n1468 & ~n1505;
  assign n1507 = ~n1467 & ~n1506;
  assign n1508 = ~n1466 & ~n1507;
  assign n1509 = ~n1465 & ~n1508;
  assign n1510 = ~n1464 & ~n1509;
  assign n1511 = ~n1463 & ~n1510;
  assign n1512 = ~n1462 & ~n1511;
  assign n1513 = ~n1461 & ~n1512;
  assign n1514 = ~n1460 & ~n1513;
  assign n1515 = ~n1459 & ~n1514;
  assign n1516 = ~n1458 & ~n1515;
  assign n1517 = ~n1457 & ~n1516;
  assign n1518 = ~n1456 & ~n1517;
  assign n1519 = ~n1455 & ~n1518;
  assign n1520 = ~n1454 & ~n1519;
  assign n1521 = ~n1453 & ~n1520;
  assign n1522 = ~n1452 & ~n1521;
  assign n1523 = ~n1451 & ~n1522;
  assign n1524 = ~n1450 & ~n1523;
  assign n1525 = ~n1449 & ~n1524;
  assign n1526 = ~n1448 & ~n1525;
  assign n1527 = ~n1447 & ~n1526;
  assign n1528 = ~n1446 & ~n1527;
  assign n1529 = ~n1445 & ~n1528;
  assign n1530 = ~n1444 & ~n1529;
  assign n1531 = ~n1442 & ~n1443;
  assign n1532 = ~n1530 & n1531;
  assign n1533 = ~n1440 & ~n1441;
  assign n1534 = ~n1532 & n1533;
  assign n1535 = pi024 & ~pi152;
  assign n1536 = pi025 & ~pi153;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = ~n1534 & n1537;
  assign n1539 = ~pi025 & pi153;
  assign n1540 = ~pi026 & pi154;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~n1538 & n1541;
  assign n1543 = pi026 & ~pi154;
  assign n1544 = pi027 & ~pi155;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = ~n1542 & n1545;
  assign n1547 = ~pi027 & pi155;
  assign n1548 = ~pi028 & pi156;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1546 & n1549;
  assign n1551 = pi028 & ~pi156;
  assign n1552 = pi029 & ~pi157;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = ~n1550 & n1553;
  assign n1555 = ~pi029 & pi157;
  assign n1556 = ~pi030 & pi158;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n1554 & n1557;
  assign n1559 = pi030 & ~pi158;
  assign n1560 = pi031 & ~pi159;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1558 & n1561;
  assign n1563 = ~pi036 & pi164;
  assign n1564 = ~pi034 & pi162;
  assign n1565 = ~pi035 & pi163;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = ~pi031 & pi159;
  assign n1568 = ~pi032 & pi160;
  assign n1569 = ~pi033 & pi161;
  assign n1570 = ~pi037 & pi165;
  assign n1571 = ~pi039 & pi167;
  assign n1572 = ~pi038 & pi166;
  assign n1573 = ~n1570 & ~n1571;
  assign n1574 = ~n1572 & n1573;
  assign n1575 = ~n1563 & ~n1567;
  assign n1576 = ~n1568 & ~n1569;
  assign n1577 = n1575 & n1576;
  assign n1578 = n1566 & n1577;
  assign n1579 = n1574 & n1578;
  assign n1580 = ~n1562 & n1579;
  assign n1581 = pi038 & ~pi166;
  assign n1582 = ~n1571 & n1581;
  assign n1583 = pi039 & ~pi167;
  assign n1584 = pi037 & ~pi165;
  assign n1585 = pi036 & ~pi164;
  assign n1586 = pi035 & ~pi163;
  assign n1587 = pi034 & ~pi162;
  assign n1588 = pi033 & ~pi161;
  assign n1589 = pi032 & ~pi160;
  assign n1590 = ~n1569 & n1589;
  assign n1591 = ~n1587 & ~n1588;
  assign n1592 = ~n1590 & n1591;
  assign n1593 = n1566 & ~n1592;
  assign n1594 = ~n1586 & ~n1593;
  assign n1595 = ~n1563 & ~n1594;
  assign n1596 = ~n1584 & ~n1585;
  assign n1597 = ~n1595 & n1596;
  assign n1598 = n1574 & ~n1597;
  assign n1599 = ~n1582 & ~n1583;
  assign n1600 = ~n1598 & n1599;
  assign n1601 = ~n1580 & n1600;
  assign n1602 = ~pi040 & pi168;
  assign n1603 = ~n1424 & ~n1602;
  assign n1604 = n1414 & n1603;
  assign n1605 = n1421 & n1604;
  assign n1606 = ~n1432 & n1605;
  assign n1607 = ~n1601 & n1606;
  assign n1608 = ~n1411 & ~n1439;
  assign n1609 = ~n1607 & n1608;
  assign n1610 = ~pi048 & pi176;
  assign n1611 = ~n1394 & ~n1610;
  assign n1612 = n1383 & n1611;
  assign n1613 = n1391 & n1612;
  assign n1614 = ~n1402 & n1613;
  assign n1615 = ~n1609 & n1614;
  assign n1616 = ~n1410 & ~n1615;
  assign n1617 = ~pi056 & pi184;
  assign n1618 = ~pi060 & pi188;
  assign n1619 = ~pi057 & pi185;
  assign n1620 = ~pi061 & pi189;
  assign n1621 = ~pi063 & pi191;
  assign n1622 = ~pi062 & pi190;
  assign n1623 = ~n1620 & ~n1621;
  assign n1624 = ~n1622 & n1623;
  assign n1625 = ~n1617 & ~n1618;
  assign n1626 = ~n1619 & n1625;
  assign n1627 = n1379 & n1626;
  assign n1628 = n1624 & n1627;
  assign n1629 = ~n1616 & n1628;
  assign n1630 = pi062 & ~pi190;
  assign n1631 = ~n1621 & n1630;
  assign n1632 = pi063 & ~pi191;
  assign n1633 = pi061 & ~pi189;
  assign n1634 = pi060 & ~pi188;
  assign n1635 = pi059 & ~pi187;
  assign n1636 = pi058 & ~pi186;
  assign n1637 = pi057 & ~pi185;
  assign n1638 = pi056 & ~pi184;
  assign n1639 = ~n1619 & n1638;
  assign n1640 = ~n1636 & ~n1637;
  assign n1641 = ~n1639 & n1640;
  assign n1642 = n1379 & ~n1641;
  assign n1643 = ~n1635 & ~n1642;
  assign n1644 = ~n1618 & ~n1643;
  assign n1645 = ~n1633 & ~n1634;
  assign n1646 = ~n1644 & n1645;
  assign n1647 = n1624 & ~n1646;
  assign n1648 = ~n1631 & ~n1632;
  assign n1649 = ~n1647 & n1648;
  assign n1650 = ~n1629 & n1649;
  assign n1651 = ~pi065 & pi193;
  assign n1652 = ~pi064 & pi192;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~n1650 & n1653;
  assign n1655 = pi066 & ~pi194;
  assign n1656 = pi065 & ~pi193;
  assign n1657 = pi064 & ~pi192;
  assign n1658 = ~n1651 & n1657;
  assign n1659 = ~n1655 & ~n1656;
  assign n1660 = ~n1658 & n1659;
  assign n1661 = ~n1654 & n1660;
  assign n1662 = ~n1376 & ~n1661;
  assign n1663 = ~n1375 & ~n1662;
  assign n1664 = ~pi069 & pi197;
  assign n1665 = ~pi068 & pi196;
  assign n1666 = ~pi070 & pi198;
  assign n1667 = ~pi071 & pi199;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~pi067 & pi195;
  assign n1670 = ~n1664 & ~n1665;
  assign n1671 = ~n1669 & n1670;
  assign n1672 = n1668 & n1671;
  assign n1673 = ~n1663 & n1672;
  assign n1674 = pi071 & ~pi199;
  assign n1675 = pi070 & ~pi198;
  assign n1676 = pi069 & ~pi197;
  assign n1677 = pi068 & ~pi196;
  assign n1678 = ~n1664 & n1677;
  assign n1679 = ~n1675 & ~n1676;
  assign n1680 = ~n1678 & n1679;
  assign n1681 = n1668 & ~n1680;
  assign n1682 = ~n1674 & ~n1681;
  assign n1683 = ~n1673 & n1682;
  assign n1684 = ~pi072 & pi200;
  assign n1685 = ~n1368 & ~n1684;
  assign n1686 = n1365 & n1685;
  assign n1687 = ~n1683 & n1686;
  assign n1688 = ~n1373 & ~n1374;
  assign n1689 = ~n1687 & n1688;
  assign n1690 = ~pi076 & pi204;
  assign n1691 = ~n1357 & ~n1690;
  assign n1692 = n1354 & n1691;
  assign n1693 = ~n1689 & n1692;
  assign n1694 = ~n1351 & ~n1362;
  assign n1695 = ~n1693 & n1694;
  assign n1696 = ~pi080 & pi208;
  assign n1697 = ~n1345 & ~n1696;
  assign n1698 = n1342 & n1697;
  assign n1699 = ~n1695 & n1698;
  assign n1700 = ~n1339 & ~n1350;
  assign n1701 = ~n1699 & n1700;
  assign n1702 = ~pi084 & pi212;
  assign n1703 = ~n1333 & ~n1702;
  assign n1704 = n1330 & n1703;
  assign n1705 = ~n1701 & n1704;
  assign n1706 = ~n1327 & ~n1338;
  assign n1707 = ~n1705 & n1706;
  assign n1708 = ~pi088 & pi216;
  assign n1709 = ~n1320 & ~n1708;
  assign n1710 = n1317 & n1709;
  assign n1711 = ~n1707 & n1710;
  assign n1712 = ~n1325 & ~n1326;
  assign n1713 = ~n1711 & n1712;
  assign n1714 = ~pi092 & pi220;
  assign n1715 = ~n1309 & ~n1714;
  assign n1716 = n1306 & n1715;
  assign n1717 = ~n1713 & n1716;
  assign n1718 = ~n1303 & ~n1314;
  assign n1719 = ~n1717 & n1718;
  assign n1720 = ~pi096 & pi224;
  assign n1721 = ~n1297 & ~n1720;
  assign n1722 = n1294 & n1721;
  assign n1723 = ~n1719 & n1722;
  assign n1724 = ~n1291 & ~n1302;
  assign n1725 = ~n1723 & n1724;
  assign n1726 = ~pi100 & pi228;
  assign n1727 = ~n1285 & ~n1726;
  assign n1728 = n1282 & n1727;
  assign n1729 = ~n1725 & n1728;
  assign n1730 = ~n1279 & ~n1290;
  assign n1731 = ~n1729 & n1730;
  assign n1732 = ~pi104 & pi232;
  assign n1733 = ~n1273 & ~n1732;
  assign n1734 = n1270 & n1733;
  assign n1735 = ~n1731 & n1734;
  assign n1736 = ~n1267 & ~n1278;
  assign n1737 = ~n1735 & n1736;
  assign n1738 = ~pi108 & pi236;
  assign n1739 = ~n1261 & ~n1738;
  assign n1740 = n1258 & n1739;
  assign n1741 = ~n1737 & n1740;
  assign n1742 = ~n1255 & ~n1266;
  assign n1743 = ~n1741 & n1742;
  assign n1744 = ~pi112 & pi240;
  assign n1745 = ~n1249 & ~n1744;
  assign n1746 = n1246 & n1745;
  assign n1747 = ~n1743 & n1746;
  assign n1748 = ~n1243 & ~n1254;
  assign n1749 = ~n1747 & n1748;
  assign n1750 = ~pi116 & pi244;
  assign n1751 = ~n1237 & ~n1750;
  assign n1752 = n1234 & n1751;
  assign n1753 = ~n1749 & n1752;
  assign n1754 = ~n1231 & ~n1242;
  assign n1755 = ~n1753 & n1754;
  assign n1756 = ~pi120 & pi248;
  assign n1757 = ~n1225 & ~n1756;
  assign n1758 = n1222 & n1757;
  assign n1759 = ~n1755 & n1758;
  assign n1760 = ~n1219 & ~n1230;
  assign n1761 = ~n1759 & n1760;
  assign n1762 = ~pi124 & pi252;
  assign n1763 = ~n1207 & ~n1762;
  assign n1764 = n1210 & n1763;
  assign n1765 = ~n1761 & n1764;
  assign n1766 = ~n1217 & ~n1218;
  assign n1767 = ~n1765 & n1766;
  assign n1768 = pi123 & ~n1767;
  assign n1769 = pi251 & n1767;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = pi379 & ~n1203;
  assign n1772 = pi507 & n1203;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = n1770 & ~n1773;
  assign n1775 = pi122 & ~n1767;
  assign n1776 = pi250 & n1767;
  assign n1777 = ~n1775 & ~n1776;
  assign n1778 = pi378 & ~n1203;
  assign n1779 = pi506 & n1203;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = n1777 & ~n1780;
  assign n1782 = ~n1774 & ~n1781;
  assign n1783 = ~n1777 & n1780;
  assign n1784 = pi121 & ~n1767;
  assign n1785 = pi249 & n1767;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = pi377 & ~n1203;
  assign n1788 = pi505 & n1203;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~n1786 & n1789;
  assign n1791 = pi376 & ~n1203;
  assign n1792 = pi504 & n1203;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = n1786 & ~n1789;
  assign n1795 = pi120 & ~n1767;
  assign n1796 = pi248 & n1767;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = n1793 & ~n1797;
  assign n1799 = ~n1794 & n1798;
  assign n1800 = ~n1783 & ~n1790;
  assign n1801 = ~n1799 & n1800;
  assign n1802 = n1782 & ~n1801;
  assign n1803 = ~n1770 & n1773;
  assign n1804 = pi119 & ~n1767;
  assign n1805 = pi247 & n1767;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = pi375 & ~n1203;
  assign n1808 = pi503 & n1203;
  assign n1809 = ~n1807 & ~n1808;
  assign n1810 = ~n1806 & n1809;
  assign n1811 = n1806 & ~n1809;
  assign n1812 = pi374 & ~n1203;
  assign n1813 = pi502 & n1203;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = pi118 & ~n1767;
  assign n1816 = pi246 & n1767;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = ~n1814 & n1817;
  assign n1819 = ~n1811 & ~n1818;
  assign n1820 = n1814 & ~n1817;
  assign n1821 = pi117 & ~n1767;
  assign n1822 = pi245 & n1767;
  assign n1823 = ~n1821 & ~n1822;
  assign n1824 = pi373 & ~n1203;
  assign n1825 = pi501 & n1203;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = ~n1823 & n1826;
  assign n1828 = pi372 & ~n1203;
  assign n1829 = pi500 & n1203;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = n1823 & ~n1826;
  assign n1832 = pi116 & ~n1767;
  assign n1833 = pi244 & n1767;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = n1830 & ~n1834;
  assign n1836 = ~n1831 & n1835;
  assign n1837 = ~n1820 & ~n1827;
  assign n1838 = ~n1836 & n1837;
  assign n1839 = n1819 & ~n1838;
  assign n1840 = pi115 & ~n1767;
  assign n1841 = pi243 & n1767;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = pi371 & ~n1203;
  assign n1844 = pi499 & n1203;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~n1842 & n1845;
  assign n1847 = n1842 & ~n1845;
  assign n1848 = pi114 & ~n1767;
  assign n1849 = pi242 & n1767;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = pi370 & ~n1203;
  assign n1852 = pi498 & n1203;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = n1850 & ~n1853;
  assign n1855 = ~n1847 & ~n1854;
  assign n1856 = ~n1850 & n1853;
  assign n1857 = pi113 & ~n1767;
  assign n1858 = pi241 & n1767;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = pi369 & ~n1203;
  assign n1861 = pi497 & n1203;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = ~n1859 & n1862;
  assign n1864 = pi368 & ~n1203;
  assign n1865 = pi496 & n1203;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = n1859 & ~n1862;
  assign n1868 = pi112 & ~n1767;
  assign n1869 = pi240 & n1767;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = n1866 & ~n1870;
  assign n1872 = ~n1867 & n1871;
  assign n1873 = ~n1856 & ~n1863;
  assign n1874 = ~n1872 & n1873;
  assign n1875 = n1855 & ~n1874;
  assign n1876 = pi107 & ~n1767;
  assign n1877 = pi235 & n1767;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = pi363 & ~n1203;
  assign n1880 = pi491 & n1203;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = n1878 & ~n1881;
  assign n1883 = pi106 & ~n1767;
  assign n1884 = pi234 & n1767;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = pi362 & ~n1203;
  assign n1887 = pi490 & n1203;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1885 & ~n1888;
  assign n1890 = ~n1882 & ~n1889;
  assign n1891 = ~n1885 & n1888;
  assign n1892 = pi105 & ~n1767;
  assign n1893 = pi233 & n1767;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = pi361 & ~n1203;
  assign n1896 = pi489 & n1203;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~n1894 & n1897;
  assign n1899 = pi360 & ~n1203;
  assign n1900 = pi488 & n1203;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = n1894 & ~n1897;
  assign n1903 = pi104 & ~n1767;
  assign n1904 = pi232 & n1767;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = n1901 & ~n1905;
  assign n1907 = ~n1902 & n1906;
  assign n1908 = ~n1891 & ~n1898;
  assign n1909 = ~n1907 & n1908;
  assign n1910 = n1890 & ~n1909;
  assign n1911 = ~n1878 & n1881;
  assign n1912 = pi103 & ~n1767;
  assign n1913 = pi231 & n1767;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = pi359 & ~n1203;
  assign n1916 = pi487 & n1203;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n1914 & n1917;
  assign n1919 = n1914 & ~n1917;
  assign n1920 = pi358 & ~n1203;
  assign n1921 = pi486 & n1203;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = pi102 & ~n1767;
  assign n1924 = pi230 & n1767;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = ~n1922 & n1925;
  assign n1927 = ~n1919 & ~n1926;
  assign n1928 = n1922 & ~n1925;
  assign n1929 = pi101 & ~n1767;
  assign n1930 = pi229 & n1767;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = pi357 & ~n1203;
  assign n1933 = pi485 & n1203;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = ~n1931 & n1934;
  assign n1936 = pi356 & ~n1203;
  assign n1937 = pi484 & n1203;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = n1931 & ~n1934;
  assign n1940 = pi100 & ~n1767;
  assign n1941 = pi228 & n1767;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = n1938 & ~n1942;
  assign n1944 = ~n1939 & n1943;
  assign n1945 = ~n1928 & ~n1935;
  assign n1946 = ~n1944 & n1945;
  assign n1947 = n1927 & ~n1946;
  assign n1948 = pi099 & ~n1767;
  assign n1949 = pi227 & n1767;
  assign n1950 = ~n1948 & ~n1949;
  assign n1951 = pi355 & ~n1203;
  assign n1952 = pi483 & n1203;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = ~n1950 & n1953;
  assign n1955 = n1950 & ~n1953;
  assign n1956 = pi098 & ~n1767;
  assign n1957 = pi226 & n1767;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = pi354 & ~n1203;
  assign n1960 = pi482 & n1203;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = n1958 & ~n1961;
  assign n1963 = ~n1955 & ~n1962;
  assign n1964 = ~n1958 & n1961;
  assign n1965 = pi097 & ~n1767;
  assign n1966 = pi225 & n1767;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = pi353 & ~n1203;
  assign n1969 = pi481 & n1203;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~n1967 & n1970;
  assign n1972 = pi352 & ~n1203;
  assign n1973 = pi480 & n1203;
  assign n1974 = ~n1972 & ~n1973;
  assign n1975 = n1967 & ~n1970;
  assign n1976 = pi096 & ~n1767;
  assign n1977 = pi224 & n1767;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = n1974 & ~n1978;
  assign n1980 = ~n1975 & n1979;
  assign n1981 = ~n1964 & ~n1971;
  assign n1982 = ~n1980 & n1981;
  assign n1983 = n1963 & ~n1982;
  assign n1984 = pi091 & ~n1767;
  assign n1985 = pi219 & n1767;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = pi347 & ~n1203;
  assign n1988 = pi475 & n1203;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = n1986 & ~n1989;
  assign n1991 = pi090 & ~n1767;
  assign n1992 = pi218 & n1767;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = pi346 & ~n1203;
  assign n1995 = pi474 & n1203;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = n1993 & ~n1996;
  assign n1998 = ~n1990 & ~n1997;
  assign n1999 = ~n1993 & n1996;
  assign n2000 = pi089 & ~n1767;
  assign n2001 = pi217 & n1767;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = pi345 & ~n1203;
  assign n2004 = pi473 & n1203;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n2002 & n2005;
  assign n2007 = pi344 & ~n1203;
  assign n2008 = pi472 & n1203;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = n2002 & ~n2005;
  assign n2011 = pi088 & ~n1767;
  assign n2012 = pi216 & n1767;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = n2009 & ~n2013;
  assign n2015 = ~n2010 & n2014;
  assign n2016 = ~n1999 & ~n2006;
  assign n2017 = ~n2015 & n2016;
  assign n2018 = n1998 & ~n2017;
  assign n2019 = ~n1986 & n1989;
  assign n2020 = pi087 & ~n1767;
  assign n2021 = pi215 & n1767;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = pi343 & ~n1203;
  assign n2024 = pi471 & n1203;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~n2022 & n2025;
  assign n2027 = n2022 & ~n2025;
  assign n2028 = pi342 & ~n1203;
  assign n2029 = pi470 & n1203;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = pi086 & ~n1767;
  assign n2032 = pi214 & n1767;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = ~n2030 & n2033;
  assign n2035 = ~n2027 & ~n2034;
  assign n2036 = n2030 & ~n2033;
  assign n2037 = pi085 & ~n1767;
  assign n2038 = pi213 & n1767;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = pi341 & ~n1203;
  assign n2041 = pi469 & n1203;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = ~n2039 & n2042;
  assign n2044 = pi340 & ~n1203;
  assign n2045 = pi468 & n1203;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = n2039 & ~n2042;
  assign n2048 = pi084 & ~n1767;
  assign n2049 = pi212 & n1767;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = n2046 & ~n2050;
  assign n2052 = ~n2047 & n2051;
  assign n2053 = ~n2036 & ~n2043;
  assign n2054 = ~n2052 & n2053;
  assign n2055 = n2035 & ~n2054;
  assign n2056 = pi083 & ~n1767;
  assign n2057 = pi211 & n1767;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = pi339 & ~n1203;
  assign n2060 = pi467 & n1203;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = ~n2058 & n2061;
  assign n2063 = n2058 & ~n2061;
  assign n2064 = pi082 & ~n1767;
  assign n2065 = pi210 & n1767;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = pi338 & ~n1203;
  assign n2068 = pi466 & n1203;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = n2066 & ~n2069;
  assign n2071 = ~n2063 & ~n2070;
  assign n2072 = ~n2066 & n2069;
  assign n2073 = pi081 & ~n1767;
  assign n2074 = pi209 & n1767;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = pi337 & ~n1203;
  assign n2077 = pi465 & n1203;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = ~n2075 & n2078;
  assign n2080 = pi336 & ~n1203;
  assign n2081 = pi464 & n1203;
  assign n2082 = ~n2080 & ~n2081;
  assign n2083 = n2075 & ~n2078;
  assign n2084 = pi080 & ~n1767;
  assign n2085 = pi208 & n1767;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = n2082 & ~n2086;
  assign n2088 = ~n2083 & n2087;
  assign n2089 = ~n2072 & ~n2079;
  assign n2090 = ~n2088 & n2089;
  assign n2091 = n2071 & ~n2090;
  assign n2092 = pi075 & ~n1767;
  assign n2093 = pi203 & n1767;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = pi331 & ~n1203;
  assign n2096 = pi459 & n1203;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = n2094 & ~n2097;
  assign n2099 = pi074 & ~n1767;
  assign n2100 = pi202 & n1767;
  assign n2101 = ~n2099 & ~n2100;
  assign n2102 = pi330 & ~n1203;
  assign n2103 = pi458 & n1203;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = n2101 & ~n2104;
  assign n2106 = ~n2098 & ~n2105;
  assign n2107 = ~n2101 & n2104;
  assign n2108 = pi073 & ~n1767;
  assign n2109 = pi201 & n1767;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = pi329 & ~n1203;
  assign n2112 = pi457 & n1203;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n2110 & n2113;
  assign n2115 = pi328 & ~n1203;
  assign n2116 = pi456 & n1203;
  assign n2117 = ~n2115 & ~n2116;
  assign n2118 = n2110 & ~n2113;
  assign n2119 = pi072 & ~n1767;
  assign n2120 = pi200 & n1767;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = n2117 & ~n2121;
  assign n2123 = ~n2118 & n2122;
  assign n2124 = ~n2107 & ~n2114;
  assign n2125 = ~n2123 & n2124;
  assign n2126 = n2106 & ~n2125;
  assign n2127 = ~n2094 & n2097;
  assign n2128 = pi067 & ~n1767;
  assign n2129 = pi195 & n1767;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = pi323 & ~n1203;
  assign n2132 = pi451 & n1203;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = n2130 & ~n2133;
  assign n2135 = pi066 & ~n1767;
  assign n2136 = pi194 & n1767;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = pi322 & ~n1203;
  assign n2139 = pi450 & n1203;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = n2137 & ~n2140;
  assign n2142 = ~n2134 & ~n2141;
  assign n2143 = ~n2137 & n2140;
  assign n2144 = pi065 & ~n1767;
  assign n2145 = pi193 & n1767;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = pi321 & ~n1203;
  assign n2148 = pi449 & n1203;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = ~n2146 & n2149;
  assign n2151 = pi320 & ~n1203;
  assign n2152 = pi448 & n1203;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = n2146 & ~n2149;
  assign n2155 = pi064 & ~n1767;
  assign n2156 = pi192 & n1767;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = n2153 & ~n2157;
  assign n2159 = ~n2154 & n2158;
  assign n2160 = ~n2143 & ~n2150;
  assign n2161 = ~n2159 & n2160;
  assign n2162 = n2142 & ~n2161;
  assign n2163 = ~n2130 & n2133;
  assign n2164 = pi285 & ~n1203;
  assign n2165 = pi413 & n1203;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = pi029 & ~n1767;
  assign n2168 = pi157 & n1767;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = n2166 & ~n2169;
  assign n2171 = pi025 & ~n1767;
  assign n2172 = pi153 & n1767;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = pi281 & ~n1203;
  assign n2175 = pi409 & n1203;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = n2173 & ~n2176;
  assign n2178 = pi024 & ~n1767;
  assign n2179 = pi152 & n1767;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = pi280 & ~n1203;
  assign n2182 = pi408 & n1203;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = ~n2180 & n2183;
  assign n2185 = pi277 & ~n1203;
  assign n2186 = pi405 & n1203;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = pi021 & ~n1767;
  assign n2189 = pi149 & n1767;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = n2187 & ~n2190;
  assign n2192 = pi017 & ~n1767;
  assign n2193 = pi145 & n1767;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = pi273 & ~n1203;
  assign n2196 = pi401 & n1203;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = n2194 & ~n2197;
  assign n2199 = pi016 & ~n1767;
  assign n2200 = pi144 & n1767;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = pi272 & ~n1203;
  assign n2203 = pi400 & n1203;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = ~n2201 & n2204;
  assign n2206 = pi269 & ~n1203;
  assign n2207 = pi397 & n1203;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = pi013 & ~n1767;
  assign n2210 = pi141 & n1767;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = n2208 & ~n2211;
  assign n2213 = pi259 & ~n1203;
  assign n2214 = pi387 & n1203;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = pi003 & ~n1767;
  assign n2217 = pi131 & n1767;
  assign n2218 = ~n2216 & ~n2217;
  assign n2219 = n2215 & ~n2218;
  assign n2220 = pi260 & ~n1203;
  assign n2221 = pi388 & n1203;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = pi004 & ~n1767;
  assign n2224 = pi132 & n1767;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = n2222 & ~n2225;
  assign n2227 = ~n2215 & n2218;
  assign n2228 = pi002 & ~n1767;
  assign n2229 = pi130 & n1767;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = pi258 & ~n1203;
  assign n2232 = pi386 & n1203;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = n2230 & ~n2233;
  assign n2235 = pi001 & ~n1767;
  assign n2236 = pi129 & n1767;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = pi257 & ~n1203;
  assign n2239 = pi385 & n1203;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = n2237 & ~n2240;
  assign n2242 = pi000 & ~n1767;
  assign n2243 = pi128 & n1767;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = n1206 & ~n2244;
  assign n2246 = ~n2241 & n2245;
  assign n2247 = ~n2230 & n2233;
  assign n2248 = ~n2237 & n2240;
  assign n2249 = ~n2247 & ~n2248;
  assign n2250 = ~n2246 & n2249;
  assign n2251 = ~n2227 & ~n2234;
  assign n2252 = ~n2250 & n2251;
  assign n2253 = ~n2219 & ~n2226;
  assign n2254 = ~n2252 & n2253;
  assign n2255 = ~n2222 & n2225;
  assign n2256 = pi005 & ~n1767;
  assign n2257 = pi133 & n1767;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = pi261 & ~n1203;
  assign n2260 = pi389 & n1203;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = n2258 & ~n2261;
  assign n2263 = ~n2255 & ~n2262;
  assign n2264 = ~n2254 & n2263;
  assign n2265 = ~n2258 & n2261;
  assign n2266 = pi262 & ~n1203;
  assign n2267 = pi390 & n1203;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = pi006 & ~n1767;
  assign n2270 = pi134 & n1767;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = n2268 & ~n2271;
  assign n2273 = ~n2265 & ~n2272;
  assign n2274 = ~n2264 & n2273;
  assign n2275 = ~n2268 & n2271;
  assign n2276 = pi263 & ~n1203;
  assign n2277 = pi391 & n1203;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = pi007 & ~n1767;
  assign n2280 = pi135 & n1767;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = ~n2278 & n2281;
  assign n2283 = ~n2275 & ~n2282;
  assign n2284 = ~n2274 & n2283;
  assign n2285 = n2278 & ~n2281;
  assign n2286 = pi008 & ~n1767;
  assign n2287 = pi136 & n1767;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = pi264 & ~n1203;
  assign n2290 = pi392 & n1203;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = ~n2288 & n2291;
  assign n2293 = ~n2285 & ~n2292;
  assign n2294 = ~n2284 & n2293;
  assign n2295 = n2288 & ~n2291;
  assign n2296 = pi009 & ~n1767;
  assign n2297 = pi137 & n1767;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = pi265 & ~n1203;
  assign n2300 = pi393 & n1203;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = n2298 & ~n2301;
  assign n2303 = ~n2295 & ~n2302;
  assign n2304 = ~n2294 & n2303;
  assign n2305 = pi010 & ~n1767;
  assign n2306 = pi138 & n1767;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = pi266 & ~n1203;
  assign n2309 = pi394 & n1203;
  assign n2310 = ~n2308 & ~n2309;
  assign n2311 = ~n2307 & n2310;
  assign n2312 = ~n2298 & n2301;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = ~n2304 & n2313;
  assign n2315 = pi267 & ~n1203;
  assign n2316 = pi395 & n1203;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = pi011 & ~n1767;
  assign n2319 = pi139 & n1767;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~n2317 & n2320;
  assign n2322 = n2307 & ~n2310;
  assign n2323 = ~n2321 & ~n2322;
  assign n2324 = ~n2314 & n2323;
  assign n2325 = n2317 & ~n2320;
  assign n2326 = pi012 & ~n1767;
  assign n2327 = pi140 & n1767;
  assign n2328 = ~n2326 & ~n2327;
  assign n2329 = pi268 & ~n1203;
  assign n2330 = pi396 & n1203;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = ~n2328 & n2331;
  assign n2333 = ~n2325 & ~n2332;
  assign n2334 = ~n2324 & n2333;
  assign n2335 = n2328 & ~n2331;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = ~n2212 & ~n2336;
  assign n2338 = ~n2208 & n2211;
  assign n2339 = pi270 & ~n1203;
  assign n2340 = pi398 & n1203;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = pi014 & ~n1767;
  assign n2343 = pi142 & n1767;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = ~n2341 & n2344;
  assign n2346 = ~n2338 & ~n2345;
  assign n2347 = ~n2337 & n2346;
  assign n2348 = n2341 & ~n2344;
  assign n2349 = pi271 & ~n1203;
  assign n2350 = pi399 & n1203;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = pi015 & ~n1767;
  assign n2353 = pi143 & n1767;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = n2351 & ~n2354;
  assign n2356 = ~n2348 & ~n2355;
  assign n2357 = ~n2347 & n2356;
  assign n2358 = ~n2351 & n2354;
  assign n2359 = n2201 & ~n2204;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~n2357 & n2360;
  assign n2362 = ~n2205 & ~n2361;
  assign n2363 = ~n2198 & ~n2362;
  assign n2364 = ~n2194 & n2197;
  assign n2365 = pi018 & ~n1767;
  assign n2366 = pi146 & n1767;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = pi274 & ~n1203;
  assign n2369 = pi402 & n1203;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = ~n2367 & n2370;
  assign n2372 = ~n2364 & ~n2371;
  assign n2373 = ~n2363 & n2372;
  assign n2374 = n2367 & ~n2370;
  assign n2375 = pi275 & ~n1203;
  assign n2376 = pi403 & n1203;
  assign n2377 = ~n2375 & ~n2376;
  assign n2378 = pi019 & ~n1767;
  assign n2379 = pi147 & n1767;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = ~n2377 & n2380;
  assign n2382 = ~n2374 & ~n2381;
  assign n2383 = ~n2373 & n2382;
  assign n2384 = n2377 & ~n2380;
  assign n2385 = pi020 & ~n1767;
  assign n2386 = pi148 & n1767;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = pi276 & ~n1203;
  assign n2389 = pi404 & n1203;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = ~n2387 & n2390;
  assign n2392 = ~n2384 & ~n2391;
  assign n2393 = ~n2383 & n2392;
  assign n2394 = n2387 & ~n2390;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = ~n2191 & ~n2395;
  assign n2397 = ~n2187 & n2190;
  assign n2398 = pi278 & ~n1203;
  assign n2399 = pi406 & n1203;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = pi022 & ~n1767;
  assign n2402 = pi150 & n1767;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~n2400 & n2403;
  assign n2405 = ~n2397 & ~n2404;
  assign n2406 = ~n2396 & n2405;
  assign n2407 = n2400 & ~n2403;
  assign n2408 = pi279 & ~n1203;
  assign n2409 = pi407 & n1203;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = pi023 & ~n1767;
  assign n2412 = pi151 & n1767;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = n2410 & ~n2413;
  assign n2415 = ~n2407 & ~n2414;
  assign n2416 = ~n2406 & n2415;
  assign n2417 = ~n2410 & n2413;
  assign n2418 = n2180 & ~n2183;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = ~n2416 & n2419;
  assign n2421 = ~n2184 & ~n2420;
  assign n2422 = ~n2177 & ~n2421;
  assign n2423 = ~n2173 & n2176;
  assign n2424 = pi026 & ~n1767;
  assign n2425 = pi154 & n1767;
  assign n2426 = ~n2424 & ~n2425;
  assign n2427 = pi282 & ~n1203;
  assign n2428 = pi410 & n1203;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n2426 & n2429;
  assign n2431 = ~n2423 & ~n2430;
  assign n2432 = ~n2422 & n2431;
  assign n2433 = n2426 & ~n2429;
  assign n2434 = pi283 & ~n1203;
  assign n2435 = pi411 & n1203;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = pi027 & ~n1767;
  assign n2438 = pi155 & n1767;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = ~n2436 & n2439;
  assign n2441 = ~n2433 & ~n2440;
  assign n2442 = ~n2432 & n2441;
  assign n2443 = n2436 & ~n2439;
  assign n2444 = pi028 & ~n1767;
  assign n2445 = pi156 & n1767;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = pi284 & ~n1203;
  assign n2448 = pi412 & n1203;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = ~n2446 & n2449;
  assign n2451 = ~n2443 & ~n2450;
  assign n2452 = ~n2442 & n2451;
  assign n2453 = n2446 & ~n2449;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = ~n2170 & ~n2454;
  assign n2456 = ~n2166 & n2169;
  assign n2457 = pi286 & ~n1203;
  assign n2458 = pi414 & n1203;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = pi030 & ~n1767;
  assign n2461 = pi158 & n1767;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = ~n2459 & n2462;
  assign n2464 = ~n2456 & ~n2463;
  assign n2465 = ~n2455 & n2464;
  assign n2466 = n2459 & ~n2462;
  assign n2467 = pi031 & ~n1767;
  assign n2468 = pi159 & n1767;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = pi287 & ~n1203;
  assign n2471 = pi415 & n1203;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = ~n2469 & n2472;
  assign n2474 = ~n2466 & ~n2473;
  assign n2475 = ~n2465 & n2474;
  assign n2476 = pi288 & ~n1203;
  assign n2477 = pi416 & n1203;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = pi032 & ~n1767;
  assign n2480 = pi160 & n1767;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = ~n2478 & n2481;
  assign n2483 = pi033 & ~n1767;
  assign n2484 = pi161 & n1767;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = pi289 & ~n1203;
  assign n2487 = pi417 & n1203;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n2485 & ~n2488;
  assign n2490 = pi035 & ~n1767;
  assign n2491 = pi163 & n1767;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = pi291 & ~n1203;
  assign n2494 = pi419 & n1203;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = n2492 & ~n2495;
  assign n2497 = pi290 & ~n1203;
  assign n2498 = pi418 & n1203;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = pi034 & ~n1767;
  assign n2501 = pi162 & n1767;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = ~n2499 & n2502;
  assign n2504 = ~n2489 & ~n2496;
  assign n2505 = ~n2503 & n2504;
  assign n2506 = pi037 & ~n1767;
  assign n2507 = pi165 & n1767;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = pi293 & ~n1203;
  assign n2510 = pi421 & n1203;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = n2508 & ~n2511;
  assign n2513 = pi039 & ~n1767;
  assign n2514 = pi167 & n1767;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = pi295 & ~n1203;
  assign n2517 = pi423 & n1203;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = n2515 & ~n2518;
  assign n2520 = pi294 & ~n1203;
  assign n2521 = pi422 & n1203;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = pi038 & ~n1767;
  assign n2524 = pi166 & n1767;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = ~n2522 & n2525;
  assign n2527 = ~n2512 & ~n2519;
  assign n2528 = ~n2526 & n2527;
  assign n2529 = n2469 & ~n2472;
  assign n2530 = pi036 & ~n1767;
  assign n2531 = pi164 & n1767;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = pi292 & ~n1203;
  assign n2534 = pi420 & n1203;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = n2532 & ~n2535;
  assign n2537 = ~n2482 & ~n2529;
  assign n2538 = ~n2536 & n2537;
  assign n2539 = n2505 & n2538;
  assign n2540 = n2528 & n2539;
  assign n2541 = ~n2475 & n2540;
  assign n2542 = n2522 & ~n2525;
  assign n2543 = ~n2519 & n2542;
  assign n2544 = ~n2515 & n2518;
  assign n2545 = ~n2532 & n2535;
  assign n2546 = ~n2508 & n2511;
  assign n2547 = n2499 & ~n2502;
  assign n2548 = ~n2496 & n2547;
  assign n2549 = ~n2492 & n2495;
  assign n2550 = n2478 & ~n2481;
  assign n2551 = ~n2485 & n2488;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = n2505 & ~n2552;
  assign n2554 = ~n2548 & ~n2549;
  assign n2555 = ~n2553 & n2554;
  assign n2556 = ~n2536 & ~n2555;
  assign n2557 = ~n2545 & ~n2546;
  assign n2558 = ~n2556 & n2557;
  assign n2559 = n2528 & ~n2558;
  assign n2560 = ~n2543 & ~n2544;
  assign n2561 = ~n2559 & n2560;
  assign n2562 = ~n2541 & n2561;
  assign n2563 = pi040 & ~n1767;
  assign n2564 = pi168 & n1767;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = pi296 & ~n1203;
  assign n2567 = pi424 & n1203;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = n2565 & ~n2568;
  assign n2570 = pi043 & ~n1767;
  assign n2571 = pi171 & n1767;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = pi299 & ~n1203;
  assign n2574 = pi427 & n1203;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = n2572 & ~n2575;
  assign n2577 = pi298 & ~n1203;
  assign n2578 = pi426 & n1203;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = pi042 & ~n1767;
  assign n2581 = pi170 & n1767;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = ~n2579 & n2582;
  assign n2584 = ~n2576 & ~n2583;
  assign n2585 = pi045 & ~n1767;
  assign n2586 = pi173 & n1767;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = pi301 & ~n1203;
  assign n2589 = pi429 & n1203;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = n2587 & ~n2590;
  assign n2592 = pi044 & ~n1767;
  assign n2593 = pi172 & n1767;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n2591 & ~n2594;
  assign n2596 = pi300 & ~n1203;
  assign n2597 = pi428 & n1203;
  assign n2598 = ~n2596 & ~n2597;
  assign n2599 = ~n2591 & n2598;
  assign n2600 = ~n2595 & ~n2599;
  assign n2601 = pi047 & ~n1767;
  assign n2602 = pi175 & n1767;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = pi303 & ~n1203;
  assign n2605 = pi431 & n1203;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n2603 & ~n2606;
  assign n2608 = pi302 & ~n1203;
  assign n2609 = pi430 & n1203;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = pi046 & ~n1767;
  assign n2612 = pi174 & n1767;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = ~n2610 & n2613;
  assign n2615 = ~n2607 & ~n2614;
  assign n2616 = pi041 & ~n1767;
  assign n2617 = pi169 & n1767;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = pi297 & ~n1203;
  assign n2620 = pi425 & n1203;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = n2618 & ~n2621;
  assign n2623 = ~n2569 & ~n2622;
  assign n2624 = n2584 & n2623;
  assign n2625 = n2615 & n2624;
  assign n2626 = ~n2600 & n2625;
  assign n2627 = ~n2562 & n2626;
  assign n2628 = ~n2603 & n2606;
  assign n2629 = n2595 & n2598;
  assign n2630 = ~n2572 & n2575;
  assign n2631 = n2579 & ~n2582;
  assign n2632 = ~n2618 & n2621;
  assign n2633 = ~n2565 & n2568;
  assign n2634 = ~n2622 & n2633;
  assign n2635 = ~n2631 & ~n2632;
  assign n2636 = ~n2634 & n2635;
  assign n2637 = n2584 & ~n2636;
  assign n2638 = ~n2630 & ~n2637;
  assign n2639 = ~n2600 & ~n2638;
  assign n2640 = n2610 & ~n2613;
  assign n2641 = ~n2587 & n2590;
  assign n2642 = ~n2640 & ~n2641;
  assign n2643 = ~n2629 & n2642;
  assign n2644 = ~n2639 & n2643;
  assign n2645 = n2615 & ~n2644;
  assign n2646 = ~n2628 & ~n2645;
  assign n2647 = ~n2627 & n2646;
  assign n2648 = pi049 & ~n1767;
  assign n2649 = pi177 & n1767;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = pi305 & ~n1203;
  assign n2652 = pi433 & n1203;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = n2650 & ~n2653;
  assign n2655 = pi051 & ~n1767;
  assign n2656 = pi179 & n1767;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = pi307 & ~n1203;
  assign n2659 = pi435 & n1203;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = n2657 & ~n2660;
  assign n2662 = pi306 & ~n1203;
  assign n2663 = pi434 & n1203;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = pi050 & ~n1767;
  assign n2666 = pi178 & n1767;
  assign n2667 = ~n2665 & ~n2666;
  assign n2668 = ~n2664 & n2667;
  assign n2669 = ~n2654 & ~n2661;
  assign n2670 = ~n2668 & n2669;
  assign n2671 = pi304 & ~n1203;
  assign n2672 = pi432 & n1203;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = pi048 & ~n1767;
  assign n2675 = pi176 & n1767;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2673 & n2676;
  assign n2678 = pi055 & ~n1767;
  assign n2679 = pi183 & n1767;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = pi311 & ~n1203;
  assign n2682 = pi439 & n1203;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = n2680 & ~n2683;
  assign n2685 = pi054 & ~n1767;
  assign n2686 = pi182 & n1767;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = pi310 & ~n1203;
  assign n2689 = pi438 & n1203;
  assign n2690 = ~n2688 & ~n2689;
  assign n2691 = n2687 & ~n2690;
  assign n2692 = ~n2684 & ~n2691;
  assign n2693 = pi053 & ~n1767;
  assign n2694 = pi181 & n1767;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = pi309 & ~n1203;
  assign n2697 = pi437 & n1203;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2695 & ~n2698;
  assign n2700 = pi308 & ~n1203;
  assign n2701 = pi436 & n1203;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = pi052 & ~n1767;
  assign n2704 = pi180 & n1767;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = ~n2702 & n2705;
  assign n2707 = ~n2699 & ~n2706;
  assign n2708 = n2692 & n2707;
  assign n2709 = n2670 & ~n2677;
  assign n2710 = n2708 & n2709;
  assign n2711 = ~n2647 & n2710;
  assign n2712 = ~n2680 & n2683;
  assign n2713 = ~n2657 & n2660;
  assign n2714 = n2673 & ~n2676;
  assign n2715 = ~n2650 & n2653;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n2670 & ~n2716;
  assign n2718 = n2664 & ~n2667;
  assign n2719 = ~n2661 & n2718;
  assign n2720 = ~n2713 & ~n2719;
  assign n2721 = ~n2717 & n2720;
  assign n2722 = n2708 & ~n2721;
  assign n2723 = ~n2687 & n2690;
  assign n2724 = ~n2695 & n2698;
  assign n2725 = n2702 & ~n2705;
  assign n2726 = ~n2699 & n2725;
  assign n2727 = ~n2723 & ~n2724;
  assign n2728 = ~n2726 & n2727;
  assign n2729 = n2692 & ~n2728;
  assign n2730 = ~n2712 & ~n2729;
  assign n2731 = ~n2722 & n2730;
  assign n2732 = ~n2711 & n2731;
  assign n2733 = pi056 & ~n1767;
  assign n2734 = pi184 & n1767;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = pi312 & ~n1203;
  assign n2737 = pi440 & n1203;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = n2735 & ~n2738;
  assign n2740 = pi059 & ~n1767;
  assign n2741 = pi187 & n1767;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = pi315 & ~n1203;
  assign n2744 = pi443 & n1203;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = n2742 & ~n2745;
  assign n2747 = pi314 & ~n1203;
  assign n2748 = pi442 & n1203;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = pi058 & ~n1767;
  assign n2751 = pi186 & n1767;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = ~n2749 & n2752;
  assign n2754 = ~n2746 & ~n2753;
  assign n2755 = pi061 & ~n1767;
  assign n2756 = pi189 & n1767;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = pi317 & ~n1203;
  assign n2759 = pi445 & n1203;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = n2757 & ~n2760;
  assign n2762 = pi060 & ~n1767;
  assign n2763 = pi188 & n1767;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = ~n2761 & ~n2764;
  assign n2766 = pi316 & ~n1203;
  assign n2767 = pi444 & n1203;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = ~n2761 & n2768;
  assign n2770 = ~n2765 & ~n2769;
  assign n2771 = pi063 & ~n1767;
  assign n2772 = pi191 & n1767;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = pi319 & ~n1203;
  assign n2775 = pi447 & n1203;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = n2773 & ~n2776;
  assign n2778 = pi318 & ~n1203;
  assign n2779 = pi446 & n1203;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = pi062 & ~n1767;
  assign n2782 = pi190 & n1767;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = ~n2780 & n2783;
  assign n2785 = ~n2777 & ~n2784;
  assign n2786 = pi057 & ~n1767;
  assign n2787 = pi185 & n1767;
  assign n2788 = ~n2786 & ~n2787;
  assign n2789 = pi313 & ~n1203;
  assign n2790 = pi441 & n1203;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = n2788 & ~n2791;
  assign n2793 = ~n2739 & ~n2792;
  assign n2794 = n2754 & n2793;
  assign n2795 = n2785 & n2794;
  assign n2796 = ~n2770 & n2795;
  assign n2797 = ~n2732 & n2796;
  assign n2798 = ~n2773 & n2776;
  assign n2799 = n2765 & n2768;
  assign n2800 = ~n2742 & n2745;
  assign n2801 = n2749 & ~n2752;
  assign n2802 = ~n2788 & n2791;
  assign n2803 = ~n2735 & n2738;
  assign n2804 = ~n2792 & n2803;
  assign n2805 = ~n2801 & ~n2802;
  assign n2806 = ~n2804 & n2805;
  assign n2807 = n2754 & ~n2806;
  assign n2808 = ~n2800 & ~n2807;
  assign n2809 = ~n2770 & ~n2808;
  assign n2810 = n2780 & ~n2783;
  assign n2811 = ~n2757 & n2760;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = ~n2799 & n2812;
  assign n2814 = ~n2809 & n2813;
  assign n2815 = n2785 & ~n2814;
  assign n2816 = ~n2798 & ~n2815;
  assign n2817 = ~n2797 & n2816;
  assign n2818 = ~n2153 & n2157;
  assign n2819 = ~n2154 & ~n2818;
  assign n2820 = n2142 & n2819;
  assign n2821 = ~n2817 & n2820;
  assign n2822 = ~n2162 & ~n2163;
  assign n2823 = ~n2821 & n2822;
  assign n2824 = pi069 & ~n1767;
  assign n2825 = pi197 & n1767;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = pi325 & ~n1203;
  assign n2828 = pi453 & n1203;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = n2826 & ~n2829;
  assign n2831 = pi068 & ~n1767;
  assign n2832 = pi196 & n1767;
  assign n2833 = ~n2831 & ~n2832;
  assign n2834 = pi324 & ~n1203;
  assign n2835 = pi452 & n1203;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = n2833 & ~n2836;
  assign n2838 = ~n2830 & ~n2837;
  assign n2839 = ~n2823 & n2838;
  assign n2840 = ~n2826 & n2829;
  assign n2841 = ~n2833 & n2836;
  assign n2842 = ~n2830 & n2841;
  assign n2843 = ~n2840 & ~n2842;
  assign n2844 = ~n2839 & n2843;
  assign n2845 = pi071 & ~n1767;
  assign n2846 = pi199 & n1767;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = pi327 & ~n1203;
  assign n2849 = pi455 & n1203;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = n2847 & ~n2850;
  assign n2852 = pi326 & ~n1203;
  assign n2853 = pi454 & n1203;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855 = pi070 & ~n1767;
  assign n2856 = pi198 & n1767;
  assign n2857 = ~n2855 & ~n2856;
  assign n2858 = ~n2854 & n2857;
  assign n2859 = ~n2851 & ~n2858;
  assign n2860 = ~n2844 & n2859;
  assign n2861 = ~n2847 & n2850;
  assign n2862 = n2854 & ~n2857;
  assign n2863 = ~n2851 & n2862;
  assign n2864 = ~n2861 & ~n2863;
  assign n2865 = ~n2860 & n2864;
  assign n2866 = ~n2117 & n2121;
  assign n2867 = ~n2118 & ~n2866;
  assign n2868 = n2106 & n2867;
  assign n2869 = ~n2865 & n2868;
  assign n2870 = ~n2126 & ~n2127;
  assign n2871 = ~n2869 & n2870;
  assign n2872 = pi077 & ~n1767;
  assign n2873 = pi205 & n1767;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = pi333 & ~n1203;
  assign n2876 = pi461 & n1203;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = n2874 & ~n2877;
  assign n2879 = pi332 & ~n1203;
  assign n2880 = pi460 & n1203;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = pi076 & ~n1767;
  assign n2883 = pi204 & n1767;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = ~n2881 & n2884;
  assign n2886 = ~n2878 & ~n2885;
  assign n2887 = ~n2871 & n2886;
  assign n2888 = ~n2874 & n2877;
  assign n2889 = n2881 & ~n2884;
  assign n2890 = ~n2878 & n2889;
  assign n2891 = ~n2888 & ~n2890;
  assign n2892 = ~n2887 & n2891;
  assign n2893 = pi079 & ~n1767;
  assign n2894 = pi207 & n1767;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = pi335 & ~n1203;
  assign n2897 = pi463 & n1203;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = n2895 & ~n2898;
  assign n2900 = pi078 & ~n1767;
  assign n2901 = pi206 & n1767;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = pi334 & ~n1203;
  assign n2904 = pi462 & n1203;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = n2902 & ~n2905;
  assign n2907 = ~n2899 & ~n2906;
  assign n2908 = ~n2892 & n2907;
  assign n2909 = ~n2895 & n2898;
  assign n2910 = ~n2902 & n2905;
  assign n2911 = ~n2899 & n2910;
  assign n2912 = ~n2909 & ~n2911;
  assign n2913 = ~n2908 & n2912;
  assign n2914 = ~n2082 & n2086;
  assign n2915 = ~n2083 & ~n2914;
  assign n2916 = n2071 & n2915;
  assign n2917 = ~n2913 & n2916;
  assign n2918 = ~n2062 & ~n2091;
  assign n2919 = ~n2917 & n2918;
  assign n2920 = ~n2046 & n2050;
  assign n2921 = ~n2047 & ~n2920;
  assign n2922 = n2035 & n2921;
  assign n2923 = ~n2919 & n2922;
  assign n2924 = ~n2026 & ~n2055;
  assign n2925 = ~n2923 & n2924;
  assign n2926 = ~n2009 & n2013;
  assign n2927 = ~n2010 & ~n2926;
  assign n2928 = n1998 & n2927;
  assign n2929 = ~n2925 & n2928;
  assign n2930 = ~n2018 & ~n2019;
  assign n2931 = ~n2929 & n2930;
  assign n2932 = pi093 & ~n1767;
  assign n2933 = pi221 & n1767;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = pi349 & ~n1203;
  assign n2936 = pi477 & n1203;
  assign n2937 = ~n2935 & ~n2936;
  assign n2938 = n2934 & ~n2937;
  assign n2939 = pi348 & ~n1203;
  assign n2940 = pi476 & n1203;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = pi092 & ~n1767;
  assign n2943 = pi220 & n1767;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n2941 & n2944;
  assign n2946 = ~n2938 & ~n2945;
  assign n2947 = ~n2931 & n2946;
  assign n2948 = ~n2934 & n2937;
  assign n2949 = n2941 & ~n2944;
  assign n2950 = ~n2938 & n2949;
  assign n2951 = ~n2948 & ~n2950;
  assign n2952 = ~n2947 & n2951;
  assign n2953 = pi095 & ~n1767;
  assign n2954 = pi223 & n1767;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = pi351 & ~n1203;
  assign n2957 = pi479 & n1203;
  assign n2958 = ~n2956 & ~n2957;
  assign n2959 = n2955 & ~n2958;
  assign n2960 = pi094 & ~n1767;
  assign n2961 = pi222 & n1767;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = pi350 & ~n1203;
  assign n2964 = pi478 & n1203;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = n2962 & ~n2965;
  assign n2967 = ~n2959 & ~n2966;
  assign n2968 = ~n2952 & n2967;
  assign n2969 = ~n2955 & n2958;
  assign n2970 = ~n2962 & n2965;
  assign n2971 = ~n2959 & n2970;
  assign n2972 = ~n2969 & ~n2971;
  assign n2973 = ~n2968 & n2972;
  assign n2974 = ~n1974 & n1978;
  assign n2975 = ~n1975 & ~n2974;
  assign n2976 = n1963 & n2975;
  assign n2977 = ~n2973 & n2976;
  assign n2978 = ~n1954 & ~n1983;
  assign n2979 = ~n2977 & n2978;
  assign n2980 = ~n1938 & n1942;
  assign n2981 = ~n1939 & ~n2980;
  assign n2982 = n1927 & n2981;
  assign n2983 = ~n2979 & n2982;
  assign n2984 = ~n1918 & ~n1947;
  assign n2985 = ~n2983 & n2984;
  assign n2986 = ~n1901 & n1905;
  assign n2987 = ~n1902 & ~n2986;
  assign n2988 = n1890 & n2987;
  assign n2989 = ~n2985 & n2988;
  assign n2990 = ~n1910 & ~n1911;
  assign n2991 = ~n2989 & n2990;
  assign n2992 = pi109 & ~n1767;
  assign n2993 = pi237 & n1767;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = pi365 & ~n1203;
  assign n2996 = pi493 & n1203;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = n2994 & ~n2997;
  assign n2999 = pi364 & ~n1203;
  assign n3000 = pi492 & n1203;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = pi108 & ~n1767;
  assign n3003 = pi236 & n1767;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = ~n3001 & n3004;
  assign n3006 = ~n2998 & ~n3005;
  assign n3007 = ~n2991 & n3006;
  assign n3008 = ~n2994 & n2997;
  assign n3009 = n3001 & ~n3004;
  assign n3010 = ~n2998 & n3009;
  assign n3011 = ~n3008 & ~n3010;
  assign n3012 = ~n3007 & n3011;
  assign n3013 = pi111 & ~n1767;
  assign n3014 = pi239 & n1767;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = pi367 & ~n1203;
  assign n3017 = pi495 & n1203;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = n3015 & ~n3018;
  assign n3020 = pi110 & ~n1767;
  assign n3021 = pi238 & n1767;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = pi366 & ~n1203;
  assign n3024 = pi494 & n1203;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = n3022 & ~n3025;
  assign n3027 = ~n3019 & ~n3026;
  assign n3028 = ~n3012 & n3027;
  assign n3029 = ~n3015 & n3018;
  assign n3030 = ~n3022 & n3025;
  assign n3031 = ~n3019 & n3030;
  assign n3032 = ~n3029 & ~n3031;
  assign n3033 = ~n3028 & n3032;
  assign n3034 = ~n1866 & n1870;
  assign n3035 = ~n1867 & ~n3034;
  assign n3036 = n1855 & n3035;
  assign n3037 = ~n3033 & n3036;
  assign n3038 = ~n1846 & ~n1875;
  assign n3039 = ~n3037 & n3038;
  assign n3040 = ~n1830 & n1834;
  assign n3041 = ~n1831 & ~n3040;
  assign n3042 = n1819 & n3041;
  assign n3043 = ~n3039 & n3042;
  assign n3044 = ~n1810 & ~n1839;
  assign n3045 = ~n3043 & n3044;
  assign n3046 = ~n1793 & n1797;
  assign n3047 = ~n1794 & ~n3046;
  assign n3048 = n1782 & n3047;
  assign n3049 = ~n3045 & n3048;
  assign n3050 = ~n1802 & ~n1803;
  assign n3051 = ~n3049 & n3050;
  assign n3052 = pi383 & pi511;
  assign n3053 = pi127 & pi255;
  assign n3054 = ~n3052 & n3053;
  assign n3055 = pi126 & ~n1767;
  assign n3056 = pi254 & n1767;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = pi382 & ~n1203;
  assign n3059 = pi510 & n1203;
  assign n3060 = ~n3058 & ~n3059;
  assign n3061 = n3057 & ~n3060;
  assign n3062 = pi381 & ~n1203;
  assign n3063 = pi509 & n1203;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = pi125 & ~n1767;
  assign n3066 = pi253 & n1767;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = ~n3064 & n3067;
  assign n3069 = ~n3061 & ~n3068;
  assign n3070 = pi124 & ~n1767;
  assign n3071 = pi252 & n1767;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = pi380 & ~n1203;
  assign n3074 = pi508 & n1203;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = n3072 & ~n3075;
  assign n3077 = ~n3054 & ~n3076;
  assign n3078 = n3069 & n3077;
  assign n3079 = ~n3051 & n3078;
  assign n3080 = n3052 & ~n3053;
  assign n3081 = ~n3072 & n3075;
  assign n3082 = n3064 & ~n3067;
  assign n3083 = ~n3081 & ~n3082;
  assign n3084 = n3069 & ~n3083;
  assign n3085 = ~n3057 & n3060;
  assign n3086 = ~n3080 & ~n3085;
  assign n3087 = ~n3084 & n3086;
  assign n3088 = ~n3054 & ~n3087;
  assign po129 = ~n3079 & ~n3088;
  assign n3090 = ~n1206 & po129;
  assign n3091 = ~n2244 & ~po129;
  assign po000 = n3090 | n3091;
  assign n3093 = ~n2240 & po129;
  assign n3094 = ~n2237 & ~po129;
  assign po001 = n3093 | n3094;
  assign n3096 = n2230 & ~po129;
  assign n3097 = n2233 & po129;
  assign po002 = ~n3096 & ~n3097;
  assign n3099 = n2218 & ~po129;
  assign n3100 = n2215 & po129;
  assign po003 = ~n3099 & ~n3100;
  assign n3102 = ~n2222 & po129;
  assign n3103 = ~n2225 & ~po129;
  assign po004 = n3102 | n3103;
  assign n3105 = ~n2261 & po129;
  assign n3106 = ~n2258 & ~po129;
  assign po005 = n3105 | n3106;
  assign n3108 = ~n2268 & po129;
  assign n3109 = ~n2271 & ~po129;
  assign po006 = n3108 | n3109;
  assign n3111 = n2281 & ~po129;
  assign n3112 = n2278 & po129;
  assign po007 = ~n3111 & ~n3112;
  assign n3114 = ~n2291 & po129;
  assign n3115 = ~n2288 & ~po129;
  assign po008 = n3114 | n3115;
  assign n3117 = n2298 & ~po129;
  assign n3118 = n2301 & po129;
  assign po009 = ~n3117 & ~n3118;
  assign n3120 = n2307 & ~po129;
  assign n3121 = n2310 & po129;
  assign po010 = ~n3120 & ~n3121;
  assign n3123 = n2320 & ~po129;
  assign n3124 = n2317 & po129;
  assign po011 = ~n3123 & ~n3124;
  assign n3126 = n2328 & ~po129;
  assign n3127 = n2331 & po129;
  assign po012 = ~n3126 & ~n3127;
  assign n3129 = n2211 & ~po129;
  assign n3130 = n2208 & po129;
  assign po013 = ~n3129 & ~n3130;
  assign n3132 = n2344 & ~po129;
  assign n3133 = n2341 & po129;
  assign po014 = ~n3132 & ~n3133;
  assign n3135 = n2354 & ~po129;
  assign n3136 = n2351 & po129;
  assign po015 = ~n3135 & ~n3136;
  assign n3138 = n2201 & ~po129;
  assign n3139 = n2204 & po129;
  assign po016 = ~n3138 & ~n3139;
  assign n3141 = n2194 & ~po129;
  assign n3142 = n2197 & po129;
  assign po017 = ~n3141 & ~n3142;
  assign n3144 = n2367 & ~po129;
  assign n3145 = n2370 & po129;
  assign po018 = ~n3144 & ~n3145;
  assign n3147 = n2380 & ~po129;
  assign n3148 = n2377 & po129;
  assign po019 = ~n3147 & ~n3148;
  assign n3150 = n2387 & ~po129;
  assign n3151 = n2390 & po129;
  assign po020 = ~n3150 & ~n3151;
  assign n3153 = n2190 & ~po129;
  assign n3154 = n2187 & po129;
  assign po021 = ~n3153 & ~n3154;
  assign n3156 = n2403 & ~po129;
  assign n3157 = n2400 & po129;
  assign po022 = ~n3156 & ~n3157;
  assign n3159 = n2413 & ~po129;
  assign n3160 = n2410 & po129;
  assign po023 = ~n3159 & ~n3160;
  assign n3162 = n2180 & ~po129;
  assign n3163 = n2183 & po129;
  assign po024 = ~n3162 & ~n3163;
  assign n3165 = n2173 & ~po129;
  assign n3166 = n2176 & po129;
  assign po025 = ~n3165 & ~n3166;
  assign n3168 = n2426 & ~po129;
  assign n3169 = n2429 & po129;
  assign po026 = ~n3168 & ~n3169;
  assign n3171 = n2439 & ~po129;
  assign n3172 = n2436 & po129;
  assign po027 = ~n3171 & ~n3172;
  assign n3174 = n2446 & ~po129;
  assign n3175 = n2449 & po129;
  assign po028 = ~n3174 & ~n3175;
  assign n3177 = n2169 & ~po129;
  assign n3178 = n2166 & po129;
  assign po029 = ~n3177 & ~n3178;
  assign n3180 = n2462 & ~po129;
  assign n3181 = n2459 & po129;
  assign po030 = ~n3180 & ~n3181;
  assign n3183 = n2469 & ~po129;
  assign n3184 = n2472 & po129;
  assign po031 = ~n3183 & ~n3184;
  assign n3186 = n2481 & ~po129;
  assign n3187 = n2478 & po129;
  assign po032 = ~n3186 & ~n3187;
  assign n3189 = n2485 & ~po129;
  assign n3190 = n2488 & po129;
  assign po033 = ~n3189 & ~n3190;
  assign n3192 = n2502 & ~po129;
  assign n3193 = n2499 & po129;
  assign po034 = ~n3192 & ~n3193;
  assign n3195 = n2492 & ~po129;
  assign n3196 = n2495 & po129;
  assign po035 = ~n3195 & ~n3196;
  assign n3198 = n2532 & ~po129;
  assign n3199 = n2535 & po129;
  assign po036 = ~n3198 & ~n3199;
  assign n3201 = n2508 & ~po129;
  assign n3202 = n2511 & po129;
  assign po037 = ~n3201 & ~n3202;
  assign n3204 = n2525 & ~po129;
  assign n3205 = n2522 & po129;
  assign po038 = ~n3204 & ~n3205;
  assign n3207 = n2515 & ~po129;
  assign n3208 = n2518 & po129;
  assign po039 = ~n3207 & ~n3208;
  assign n3210 = n2565 & ~po129;
  assign n3211 = n2568 & po129;
  assign po040 = ~n3210 & ~n3211;
  assign n3213 = n2618 & ~po129;
  assign n3214 = n2621 & po129;
  assign po041 = ~n3213 & ~n3214;
  assign n3216 = n2582 & ~po129;
  assign n3217 = n2579 & po129;
  assign po042 = ~n3216 & ~n3217;
  assign n3219 = n2572 & ~po129;
  assign n3220 = n2575 & po129;
  assign po043 = ~n3219 & ~n3220;
  assign n3222 = n2594 & ~po129;
  assign n3223 = n2598 & po129;
  assign po044 = ~n3222 & ~n3223;
  assign n3225 = n2587 & ~po129;
  assign n3226 = n2590 & po129;
  assign po045 = ~n3225 & ~n3226;
  assign n3228 = n2613 & ~po129;
  assign n3229 = n2610 & po129;
  assign po046 = ~n3228 & ~n3229;
  assign n3231 = n2603 & ~po129;
  assign n3232 = n2606 & po129;
  assign po047 = ~n3231 & ~n3232;
  assign n3234 = n2676 & ~po129;
  assign n3235 = n2673 & po129;
  assign po048 = ~n3234 & ~n3235;
  assign n3237 = n2650 & ~po129;
  assign n3238 = n2653 & po129;
  assign po049 = ~n3237 & ~n3238;
  assign n3240 = n2667 & ~po129;
  assign n3241 = n2664 & po129;
  assign po050 = ~n3240 & ~n3241;
  assign n3243 = n2657 & ~po129;
  assign n3244 = n2660 & po129;
  assign po051 = ~n3243 & ~n3244;
  assign n3246 = n2705 & ~po129;
  assign n3247 = n2702 & po129;
  assign po052 = ~n3246 & ~n3247;
  assign n3249 = n2695 & ~po129;
  assign n3250 = n2698 & po129;
  assign po053 = ~n3249 & ~n3250;
  assign n3252 = n2687 & ~po129;
  assign n3253 = n2690 & po129;
  assign po054 = ~n3252 & ~n3253;
  assign n3255 = n2680 & ~po129;
  assign n3256 = n2683 & po129;
  assign po055 = ~n3255 & ~n3256;
  assign n3258 = n2735 & ~po129;
  assign n3259 = n2738 & po129;
  assign po056 = ~n3258 & ~n3259;
  assign n3261 = n2788 & ~po129;
  assign n3262 = n2791 & po129;
  assign po057 = ~n3261 & ~n3262;
  assign n3264 = n2752 & ~po129;
  assign n3265 = n2749 & po129;
  assign po058 = ~n3264 & ~n3265;
  assign n3267 = n2742 & ~po129;
  assign n3268 = n2745 & po129;
  assign po059 = ~n3267 & ~n3268;
  assign n3270 = n2764 & ~po129;
  assign n3271 = n2768 & po129;
  assign po060 = ~n3270 & ~n3271;
  assign n3273 = n2757 & ~po129;
  assign n3274 = n2760 & po129;
  assign po061 = ~n3273 & ~n3274;
  assign n3276 = n2783 & ~po129;
  assign n3277 = n2780 & po129;
  assign po062 = ~n3276 & ~n3277;
  assign n3279 = n2773 & ~po129;
  assign n3280 = n2776 & po129;
  assign po063 = ~n3279 & ~n3280;
  assign n3282 = n2157 & ~po129;
  assign n3283 = n2153 & po129;
  assign po064 = ~n3282 & ~n3283;
  assign n3285 = n2146 & ~po129;
  assign n3286 = n2149 & po129;
  assign po065 = ~n3285 & ~n3286;
  assign n3288 = n2137 & ~po129;
  assign n3289 = n2140 & po129;
  assign po066 = ~n3288 & ~n3289;
  assign n3291 = n2130 & ~po129;
  assign n3292 = n2133 & po129;
  assign po067 = ~n3291 & ~n3292;
  assign n3294 = n2833 & ~po129;
  assign n3295 = n2836 & po129;
  assign po068 = ~n3294 & ~n3295;
  assign n3297 = n2826 & ~po129;
  assign n3298 = n2829 & po129;
  assign po069 = ~n3297 & ~n3298;
  assign n3300 = n2857 & ~po129;
  assign n3301 = n2854 & po129;
  assign po070 = ~n3300 & ~n3301;
  assign n3303 = n2847 & ~po129;
  assign n3304 = n2850 & po129;
  assign po071 = ~n3303 & ~n3304;
  assign n3306 = n2121 & ~po129;
  assign n3307 = n2117 & po129;
  assign po072 = ~n3306 & ~n3307;
  assign n3309 = n2110 & ~po129;
  assign n3310 = n2113 & po129;
  assign po073 = ~n3309 & ~n3310;
  assign n3312 = n2101 & ~po129;
  assign n3313 = n2104 & po129;
  assign po074 = ~n3312 & ~n3313;
  assign n3315 = n2094 & ~po129;
  assign n3316 = n2097 & po129;
  assign po075 = ~n3315 & ~n3316;
  assign n3318 = n2884 & ~po129;
  assign n3319 = n2881 & po129;
  assign po076 = ~n3318 & ~n3319;
  assign n3321 = n2874 & ~po129;
  assign n3322 = n2877 & po129;
  assign po077 = ~n3321 & ~n3322;
  assign n3324 = n2902 & ~po129;
  assign n3325 = n2905 & po129;
  assign po078 = ~n3324 & ~n3325;
  assign n3327 = n2895 & ~po129;
  assign n3328 = n2898 & po129;
  assign po079 = ~n3327 & ~n3328;
  assign n3330 = n2086 & ~po129;
  assign n3331 = n2082 & po129;
  assign po080 = ~n3330 & ~n3331;
  assign n3333 = n2075 & ~po129;
  assign n3334 = n2078 & po129;
  assign po081 = ~n3333 & ~n3334;
  assign n3336 = n2066 & ~po129;
  assign n3337 = n2069 & po129;
  assign po082 = ~n3336 & ~n3337;
  assign n3339 = n2058 & ~po129;
  assign n3340 = n2061 & po129;
  assign po083 = ~n3339 & ~n3340;
  assign n3342 = n2050 & ~po129;
  assign n3343 = n2046 & po129;
  assign po084 = ~n3342 & ~n3343;
  assign n3345 = n2039 & ~po129;
  assign n3346 = n2042 & po129;
  assign po085 = ~n3345 & ~n3346;
  assign n3348 = n2033 & ~po129;
  assign n3349 = n2030 & po129;
  assign po086 = ~n3348 & ~n3349;
  assign n3351 = n2022 & ~po129;
  assign n3352 = n2025 & po129;
  assign po087 = ~n3351 & ~n3352;
  assign n3354 = n2013 & ~po129;
  assign n3355 = n2009 & po129;
  assign po088 = ~n3354 & ~n3355;
  assign n3357 = n2002 & ~po129;
  assign n3358 = n2005 & po129;
  assign po089 = ~n3357 & ~n3358;
  assign n3360 = n1993 & ~po129;
  assign n3361 = n1996 & po129;
  assign po090 = ~n3360 & ~n3361;
  assign n3363 = n1986 & ~po129;
  assign n3364 = n1989 & po129;
  assign po091 = ~n3363 & ~n3364;
  assign n3366 = n2944 & ~po129;
  assign n3367 = n2941 & po129;
  assign po092 = ~n3366 & ~n3367;
  assign n3369 = n2934 & ~po129;
  assign n3370 = n2937 & po129;
  assign po093 = ~n3369 & ~n3370;
  assign n3372 = n2962 & ~po129;
  assign n3373 = n2965 & po129;
  assign po094 = ~n3372 & ~n3373;
  assign n3375 = n2955 & ~po129;
  assign n3376 = n2958 & po129;
  assign po095 = ~n3375 & ~n3376;
  assign n3378 = n1978 & ~po129;
  assign n3379 = n1974 & po129;
  assign po096 = ~n3378 & ~n3379;
  assign n3381 = n1967 & ~po129;
  assign n3382 = n1970 & po129;
  assign po097 = ~n3381 & ~n3382;
  assign n3384 = n1958 & ~po129;
  assign n3385 = n1961 & po129;
  assign po098 = ~n3384 & ~n3385;
  assign n3387 = n1950 & ~po129;
  assign n3388 = n1953 & po129;
  assign po099 = ~n3387 & ~n3388;
  assign n3390 = n1942 & ~po129;
  assign n3391 = n1938 & po129;
  assign po100 = ~n3390 & ~n3391;
  assign n3393 = n1931 & ~po129;
  assign n3394 = n1934 & po129;
  assign po101 = ~n3393 & ~n3394;
  assign n3396 = n1925 & ~po129;
  assign n3397 = n1922 & po129;
  assign po102 = ~n3396 & ~n3397;
  assign n3399 = n1914 & ~po129;
  assign n3400 = n1917 & po129;
  assign po103 = ~n3399 & ~n3400;
  assign n3402 = n1905 & ~po129;
  assign n3403 = n1901 & po129;
  assign po104 = ~n3402 & ~n3403;
  assign n3405 = n1894 & ~po129;
  assign n3406 = n1897 & po129;
  assign po105 = ~n3405 & ~n3406;
  assign n3408 = n1885 & ~po129;
  assign n3409 = n1888 & po129;
  assign po106 = ~n3408 & ~n3409;
  assign n3411 = n1878 & ~po129;
  assign n3412 = n1881 & po129;
  assign po107 = ~n3411 & ~n3412;
  assign n3414 = n3004 & ~po129;
  assign n3415 = n3001 & po129;
  assign po108 = ~n3414 & ~n3415;
  assign n3417 = n2994 & ~po129;
  assign n3418 = n2997 & po129;
  assign po109 = ~n3417 & ~n3418;
  assign n3420 = n3022 & ~po129;
  assign n3421 = n3025 & po129;
  assign po110 = ~n3420 & ~n3421;
  assign n3423 = n3015 & ~po129;
  assign n3424 = n3018 & po129;
  assign po111 = ~n3423 & ~n3424;
  assign n3426 = n1870 & ~po129;
  assign n3427 = n1866 & po129;
  assign po112 = ~n3426 & ~n3427;
  assign n3429 = n1859 & ~po129;
  assign n3430 = n1862 & po129;
  assign po113 = ~n3429 & ~n3430;
  assign n3432 = n1850 & ~po129;
  assign n3433 = n1853 & po129;
  assign po114 = ~n3432 & ~n3433;
  assign n3435 = n1842 & ~po129;
  assign n3436 = n1845 & po129;
  assign po115 = ~n3435 & ~n3436;
  assign n3438 = n1834 & ~po129;
  assign n3439 = n1830 & po129;
  assign po116 = ~n3438 & ~n3439;
  assign n3441 = n1823 & ~po129;
  assign n3442 = n1826 & po129;
  assign po117 = ~n3441 & ~n3442;
  assign n3444 = n1817 & ~po129;
  assign n3445 = n1814 & po129;
  assign po118 = ~n3444 & ~n3445;
  assign n3447 = n1806 & ~po129;
  assign n3448 = n1809 & po129;
  assign po119 = ~n3447 & ~n3448;
  assign n3450 = n1797 & ~po129;
  assign n3451 = n1793 & po129;
  assign po120 = ~n3450 & ~n3451;
  assign n3453 = n1786 & ~po129;
  assign n3454 = n1789 & po129;
  assign po121 = ~n3453 & ~n3454;
  assign n3456 = n1777 & ~po129;
  assign n3457 = n1780 & po129;
  assign po122 = ~n3456 & ~n3457;
  assign n3459 = n1770 & ~po129;
  assign n3460 = n1773 & po129;
  assign po123 = ~n3459 & ~n3460;
  assign n3462 = n3072 & ~po129;
  assign n3463 = n3075 & po129;
  assign po124 = ~n3462 & ~n3463;
  assign n3465 = n3067 & ~po129;
  assign n3466 = n3064 & po129;
  assign po125 = ~n3465 & ~n3466;
  assign n3468 = n3057 & ~po129;
  assign n3469 = n3060 & po129;
  assign po126 = ~n3468 & ~n3469;
  assign po127 = n3052 & n3053;
  assign n3472 = n1767 & ~po129;
  assign n3473 = n1203 & po129;
  assign po128 = n3472 | n3473;
endmodule


