// Benchmark "y0" written by ABC on Wed Apr 26 16:30:55 2017

module y0 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159;
  wire n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1126, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
    n1553, n1554, n1555, n1556, n1557, n1558, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1821, n1822, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2222, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2464, n2465, n2466,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2484, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
    n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
    n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
    n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
    n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
    n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
    n3702, n3703, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
    n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
    n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
    n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
    n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
    n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
    n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
    n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
    n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
    n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
    n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
    n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
    n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
    n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
    n4535, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
    n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
    n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
    n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
    n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
    n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
    n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5152, n5153, n5154, n5155, n5156, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
    n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
    n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
    n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
    n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
    n5355, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
    n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5968, n5969,
    n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
    n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6120, n6121, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
    n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
    n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
    n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
    n6359, n6360, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
    n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
    n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
    n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
    n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
    n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
    n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
    n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
    n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
    n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
    n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
    n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6799, n6800, n6801, n6802, n6803,
    n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829, n6831, n6832, n6833, n6834,
    n6835, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852, n6854, n6855, n6856, n6858,
    n6859, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
    n6870, n6871, n6873, n6874, n6875, n6876, n6878, n6879, n6880, n6881,
    n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
    n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
    n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
    n6943, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
    n6954, n6955, n6956, n6957, n6959, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7115, n7116, n7119, n7120, n7121, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
    n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7262, n7263, n7264, n7265, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
    n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
    n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
    n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7388, n7389, n7390, n7391, n7392, n7394, n7395,
    n7398, n7399, n7400, n7402, n7404, n7405, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7424, n7425, n7426, n7428, n7429, n7430, n7431,
    n7432, n7434, n7435, n7437, n7438, n7440, n7441, n7442, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7480, n7481, n7482, n7483, n7484, n7485, n7487, n7488, n7489,
    n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
    n7500, n7501, n7502, n7503, n7504, n7506, n7508, n7509, n7510, n7511,
    n7512, n7513, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7551, n7552, n7553,
    n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
    n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
    n7644, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
    n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
    n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7833, n7834, n7835,
    n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
    n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
    n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
    n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
    n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
    n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
    n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8028, n8029, n8030, n8031, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
    n8048, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
    n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
    n8293, n8294, n8295, n8296, n8298, n8299, n8300, n8301, n8302, n8303,
    n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8325,
    n8326, n8327, n8328, n8329, n8331, n8332, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8346, n8347, n8348,
    n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8404, n8405, n8406, n8407, n8409, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8424;
  assign n290 = pi009 & ~pi010;
  assign n291 = ~pi007 & n290;
  assign n292 = ~pi005 & pi006;
  assign n293 = ~pi004 & n292;
  assign n294 = pi000 & pi002;
  assign n295 = pi003 & ~pi127;
  assign n296 = n294 & n295;
  assign n297 = ~pi001 & n296;
  assign n298 = n293 & n297;
  assign n299 = ~pi008 & n298;
  assign n300 = pi014 & n299;
  assign n301 = n291 & n300;
  assign n302 = ~pi012 & ~pi013;
  assign n303 = pi011 & ~pi015;
  assign n304 = n302 & n303;
  assign n305 = n301 & n304;
  assign n306 = pi001 & ~pi007;
  assign n307 = pi005 & ~pi006;
  assign n308 = ~pi004 & n307;
  assign n309 = ~pi000 & ~pi127;
  assign n310 = ~pi002 & n309;
  assign n311 = ~pi003 & n310;
  assign n312 = n308 & n311;
  assign n313 = n306 & n312;
  assign n314 = ~pi004 & pi005;
  assign n315 = pi006 & n314;
  assign n316 = pi000 & ~pi127;
  assign n317 = ~pi002 & n316;
  assign n318 = ~pi003 & n306;
  assign n319 = n317 & n318;
  assign n320 = n315 & n319;
  assign n321 = ~pi014 & ~pi015;
  assign n322 = n302 & n321;
  assign n323 = n320 & n322;
  assign n324 = ~n313 & ~n323;
  assign n325 = ~pi031 & ~n324;
  assign n326 = ~pi024 & ~pi028;
  assign n327 = ~pi025 & ~pi026;
  assign n328 = n326 & n327;
  assign n329 = ~pi027 & n328;
  assign n330 = pi029 & n329;
  assign n331 = n325 & n330;
  assign n332 = pi012 & pi013;
  assign n333 = pi002 & n316;
  assign n334 = ~pi003 & n333;
  assign n335 = ~pi001 & pi007;
  assign n336 = ~pi004 & pi006;
  assign n337 = n335 & n336;
  assign n338 = pi005 & n337;
  assign n339 = n334 & n338;
  assign n340 = ~pi014 & n339;
  assign n341 = n332 & n340;
  assign n342 = ~n331 & ~n341;
  assign n343 = ~n305 & n342;
  assign n344 = pi044 & pi045;
  assign n345 = pi122 & ~n344;
  assign n346 = n293 & n345;
  assign n347 = pi021 & ~pi022;
  assign n348 = ~pi023 & n347;
  assign n349 = pi001 & pi007;
  assign n350 = ~pi003 & n349;
  assign n351 = n333 & n350;
  assign n352 = ~pi016 & n351;
  assign n353 = pi019 & n352;
  assign n354 = pi017 & n353;
  assign n355 = pi020 & n354;
  assign n356 = n348 & n355;
  assign n357 = pi018 & n356;
  assign n358 = n346 & n357;
  assign n359 = ~pi018 & pi020;
  assign n360 = pi122 & n344;
  assign n361 = n293 & ~n360;
  assign n362 = ~pi017 & n352;
  assign n363 = n361 & n362;
  assign n364 = n348 & n363;
  assign n365 = n359 & n364;
  assign n366 = ~n358 & ~n365;
  assign n367 = n343 & n366;
  assign n368 = pi015 & n332;
  assign n369 = ~pi001 & ~pi007;
  assign n370 = n315 & n369;
  assign n371 = n334 & n370;
  assign n372 = pi014 & n371;
  assign n373 = n345 & n372;
  assign n374 = n368 & n373;
  assign n375 = ~pi003 & n309;
  assign n376 = pi004 & n307;
  assign n377 = n306 & n376;
  assign n378 = n375 & n377;
  assign n379 = n345 & n378;
  assign n380 = ~pi002 & n379;
  assign n381 = pi044 & ~pi122;
  assign n382 = ~pi018 & n356;
  assign n383 = n293 & n382;
  assign n384 = ~pi018 & pi022;
  assign n385 = ~pi020 & pi021;
  assign n386 = n384 & n385;
  assign n387 = n293 & n386;
  assign n388 = ~pi023 & n387;
  assign n389 = ~pi017 & n351;
  assign n390 = pi016 & n389;
  assign n391 = n388 & n390;
  assign n392 = n310 & n377;
  assign n393 = pi003 & n392;
  assign n394 = ~n391 & ~n393;
  assign n395 = ~n383 & n394;
  assign n396 = ~n381 & ~n395;
  assign n397 = ~pi122 & n392;
  assign n398 = ~n380 & ~n397;
  assign n399 = ~n396 & n398;
  assign n400 = pi016 & pi023;
  assign n401 = n389 & n400;
  assign n402 = n387 & n401;
  assign n403 = n349 & n376;
  assign n404 = pi003 & n309;
  assign n405 = ~pi002 & n404;
  assign n406 = n403 & n405;
  assign n407 = ~n402 & ~n406;
  assign n408 = pi027 & n328;
  assign n409 = ~n407 & n408;
  assign n410 = n347 & n359;
  assign n411 = n362 & n410;
  assign n412 = pi023 & n411;
  assign n413 = n293 & n412;
  assign n414 = n408 & n413;
  assign n415 = ~n409 & ~n414;
  assign n416 = pi004 & n292;
  assign n417 = pi021 & n359;
  assign n418 = pi017 & n351;
  assign n419 = pi016 & n418;
  assign n420 = pi019 & n419;
  assign n421 = n417 & n420;
  assign n422 = ~n411 & ~n421;
  assign n423 = n416 & ~n422;
  assign n424 = n415 & ~n423;
  assign n425 = n318 & n333;
  assign n426 = pi017 & n425;
  assign n427 = pi019 & n376;
  assign n428 = ~pi016 & n427;
  assign n429 = n426 & n428;
  assign n430 = ~pi018 & n429;
  assign n431 = ~pi022 & pi023;
  assign n432 = n430 & n431;
  assign n433 = n424 & ~n432;
  assign n434 = pi022 & n359;
  assign n435 = pi023 & n434;
  assign n436 = n363 & n435;
  assign n437 = pi008 & n298;
  assign n438 = pi014 & n437;
  assign n439 = n291 & n438;
  assign n440 = n368 & n439;
  assign n441 = ~pi011 & n440;
  assign n442 = pi012 & ~pi013;
  assign n443 = pi014 & n319;
  assign n444 = pi015 & n443;
  assign n445 = n307 & n442;
  assign n446 = n444 & n445;
  assign n447 = pi004 & n446;
  assign n448 = pi011 & ~pi013;
  assign n449 = ~pi012 & pi015;
  assign n450 = n448 & n449;
  assign n451 = n329 & n450;
  assign n452 = pi003 & n335;
  assign n453 = ~pi005 & ~pi006;
  assign n454 = pi004 & n453;
  assign n455 = n452 & n454;
  assign n456 = n333 & n455;
  assign n457 = ~pi008 & n456;
  assign n458 = pi014 & n457;
  assign n459 = ~pi010 & n458;
  assign n460 = ~pi009 & n459;
  assign n461 = n451 & n460;
  assign n462 = ~n441 & ~n447;
  assign n463 = ~n461 & n462;
  assign n464 = pi011 & n302;
  assign n465 = ~pi009 & ~pi010;
  assign n466 = n457 & n465;
  assign n467 = ~pi014 & n466;
  assign n468 = n464 & n467;
  assign n469 = n385 & ~n431;
  assign n470 = n430 & n469;
  assign n471 = ~n468 & ~n470;
  assign n472 = n329 & ~n471;
  assign n473 = pi045 & pi122;
  assign n474 = pi044 & n473;
  assign n475 = pi003 & n306;
  assign n476 = n310 & n475;
  assign n477 = pi007 & n297;
  assign n478 = ~n476 & ~n477;
  assign n479 = pi004 & pi005;
  assign n480 = pi006 & n479;
  assign n481 = ~n478 & n480;
  assign n482 = pi021 & pi022;
  assign n483 = n293 & n482;
  assign n484 = ~pi018 & n483;
  assign n485 = pi019 & pi023;
  assign n486 = n418 & n485;
  assign n487 = ~pi016 & n486;
  assign n488 = n484 & n487;
  assign n489 = ~n481 & ~n488;
  assign n490 = ~n474 & ~n489;
  assign n491 = ~pi027 & ~pi029;
  assign n492 = n328 & n491;
  assign n493 = ~pi012 & pi013;
  assign n494 = ~pi015 & n493;
  assign n495 = n376 & n494;
  assign n496 = n443 & n495;
  assign n497 = n492 & n496;
  assign n498 = ~pi039 & n311;
  assign n499 = ~pi007 & n498;
  assign n500 = pi039 & n311;
  assign n501 = n306 & n500;
  assign n502 = ~n499 & ~n501;
  assign n503 = n315 & n492;
  assign n504 = ~n502 & n503;
  assign n505 = ~n497 & ~n504;
  assign n506 = n354 & n361;
  assign n507 = ~pi018 & ~pi020;
  assign n508 = pi021 & n507;
  assign n509 = ~pi023 & n508;
  assign n510 = ~pi021 & pi022;
  assign n511 = n359 & n510;
  assign n512 = ~n509 & ~n511;
  assign n513 = n506 & ~n512;
  assign n514 = ~pi023 & n353;
  assign n515 = n359 & n483;
  assign n516 = ~n360 & n515;
  assign n517 = n514 & n516;
  assign n518 = pi004 & ~pi005;
  assign n519 = ~pi003 & n317;
  assign n520 = ~pi001 & n519;
  assign n521 = n369 & n405;
  assign n522 = ~n520 & ~n521;
  assign n523 = n518 & ~n522;
  assign n524 = ~n314 & ~n518;
  assign n525 = n310 & n452;
  assign n526 = pi006 & ~n524;
  assign n527 = n525 & n526;
  assign n528 = n314 & n405;
  assign n529 = n306 & ~n474;
  assign n530 = ~n369 & ~n529;
  assign n531 = n528 & ~n530;
  assign n532 = pi125 & ~pi126;
  assign n533 = ~pi125 & pi126;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~pi025 & n326;
  assign n536 = pi026 & ~pi027;
  assign n537 = n535 & n536;
  assign n538 = ~n534 & n537;
  assign n539 = ~n527 & ~n538;
  assign n540 = ~n531 & n539;
  assign n541 = ~n523 & n540;
  assign n542 = ~n436 & n541;
  assign n543 = ~n517 & n542;
  assign n544 = n505 & ~n513;
  assign n545 = n543 & n544;
  assign n546 = ~n490 & n545;
  assign n547 = ~n472 & n546;
  assign n548 = n463 & n547;
  assign n549 = ~pi004 & n453;
  assign n550 = pi002 & n404;
  assign n551 = n349 & ~n474;
  assign n552 = n550 & n551;
  assign n553 = n549 & n552;
  assign n554 = ~pi001 & n404;
  assign n555 = ~pi002 & n554;
  assign n556 = n524 & n555;
  assign n557 = pi019 & n391;
  assign n558 = ~pi122 & n557;
  assign n559 = ~n553 & ~n556;
  assign n560 = ~n374 & n559;
  assign n561 = ~n558 & n560;
  assign n562 = n367 & n561;
  assign n563 = n433 & n562;
  assign n564 = n399 & n548;
  assign n565 = n563 & n564;
  assign n566 = pi018 & ~pi020;
  assign n567 = ~pi021 & ~pi022;
  assign n568 = n566 & n567;
  assign n569 = n362 & n568;
  assign n570 = n485 & n569;
  assign n571 = ~n477 & ~n570;
  assign n572 = n329 & n416;
  assign n573 = pi029 & n572;
  assign n574 = ~n571 & n573;
  assign n575 = ~pi021 & n359;
  assign n576 = pi016 & n426;
  assign n577 = n427 & n576;
  assign n578 = n575 & n577;
  assign n579 = pi014 & n465;
  assign n580 = ~pi011 & ~pi015;
  assign n581 = n302 & n580;
  assign n582 = n579 & n581;
  assign n583 = n456 & n582;
  assign n584 = ~pi011 & pi015;
  assign n585 = n442 & n584;
  assign n586 = n467 & n585;
  assign n587 = ~n583 & ~n586;
  assign n588 = ~n578 & n587;
  assign n589 = ~pi015 & n442;
  assign n590 = n319 & n589;
  assign n591 = n376 & n590;
  assign n592 = ~pi019 & n362;
  assign n593 = n416 & n592;
  assign n594 = n511 & n593;
  assign n595 = ~n591 & ~n594;
  assign n596 = n347 & n507;
  assign n597 = ~n568 & ~n596;
  assign n598 = pi019 & ~pi023;
  assign n599 = n362 & n598;
  assign n600 = ~n597 & n599;
  assign n601 = ~pi007 & n297;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~pi029 & n572;
  assign n604 = ~n360 & n603;
  assign n605 = ~n602 & n604;
  assign n606 = ~pi011 & n493;
  assign n607 = ~pi009 & pi010;
  assign n608 = n606 & n607;
  assign n609 = ~pi014 & n299;
  assign n610 = ~pi015 & n608;
  assign n611 = n609 & n610;
  assign n612 = ~pi007 & n611;
  assign n613 = ~n605 & ~n612;
  assign n614 = n595 & n613;
  assign n615 = ~pi023 & n363;
  assign n616 = ~pi018 & n510;
  assign n617 = n615 & n616;
  assign n618 = n588 & ~n617;
  assign n619 = n614 & n618;
  assign n620 = pi008 & n456;
  assign n621 = pi009 & n620;
  assign n622 = ~pi010 & n621;
  assign n623 = ~n339 & ~n622;
  assign n624 = n442 & ~n623;
  assign n625 = ~pi011 & n302;
  assign n626 = ~n585 & ~n625;
  assign n627 = n291 & n437;
  assign n628 = ~pi014 & n627;
  assign n629 = ~n626 & n628;
  assign n630 = n359 & n567;
  assign n631 = n363 & n630;
  assign n632 = n310 & n416;
  assign n633 = n306 & n632;
  assign n634 = ~n474 & n633;
  assign n635 = ~n631 & ~n634;
  assign n636 = pi016 & ~pi019;
  assign n637 = n376 & n636;
  assign n638 = ~pi021 & n507;
  assign n639 = n637 & n638;
  assign n640 = n418 & n639;
  assign n641 = n345 & n640;
  assign n642 = pi022 & ~pi023;
  assign n643 = n507 & n642;
  assign n644 = n389 & n636;
  assign n645 = n643 & n644;
  assign n646 = ~pi122 & n293;
  assign n647 = ~pi021 & n346;
  assign n648 = ~n646 & ~n647;
  assign n649 = n645 & ~n648;
  assign n650 = ~n641 & ~n649;
  assign n651 = n635 & n650;
  assign n652 = ~pi012 & n303;
  assign n653 = pi011 & pi015;
  assign n654 = pi013 & n653;
  assign n655 = ~n584 & ~n652;
  assign n656 = ~n654 & n655;
  assign n657 = n465 & ~n656;
  assign n658 = ~n608 & ~n657;
  assign n659 = n458 & ~n658;
  assign n660 = ~n442 & ~n606;
  assign n661 = ~n584 & ~n660;
  assign n662 = n466 & n661;
  assign n663 = ~n659 & ~n662;
  assign n664 = ~pi014 & n620;
  assign n665 = n465 & n664;
  assign n666 = n493 & n665;
  assign n667 = pi018 & pi020;
  assign n668 = ~pi021 & n667;
  assign n669 = ~pi023 & n668;
  assign n670 = n506 & n669;
  assign n671 = pi022 & n670;
  assign n672 = pi015 & n493;
  assign n673 = n442 & ~n580;
  assign n674 = ~n672 & ~n673;
  assign n675 = pi009 & pi010;
  assign n676 = pi008 & n675;
  assign n677 = n456 & n676;
  assign n678 = pi014 & n677;
  assign n679 = ~n674 & n678;
  assign n680 = pi011 & ~pi012;
  assign n681 = ~pi013 & ~n680;
  assign n682 = ~pi014 & n456;
  assign n683 = n676 & n682;
  assign n684 = n681 & n683;
  assign n685 = ~n580 & n684;
  assign n686 = ~n679 & ~n685;
  assign n687 = ~pi004 & ~pi005;
  assign n688 = n442 & n687;
  assign n689 = n319 & n688;
  assign n690 = pi006 & n689;
  assign n691 = n686 & ~n690;
  assign n692 = ~pi011 & n442;
  assign n693 = ~pi015 & n692;
  assign n694 = ~n494 & ~n693;
  assign n695 = n677 & ~n694;
  assign n696 = n691 & ~n695;
  assign n697 = n356 & n646;
  assign n698 = pi023 & n506;
  assign n699 = pi018 & n510;
  assign n700 = n698 & n699;
  assign n701 = ~n697 & ~n700;
  assign n702 = ~pi011 & n332;
  assign n703 = pi011 & pi013;
  assign n704 = ~n449 & n703;
  assign n705 = ~n702 & ~n704;
  assign n706 = n467 & ~n705;
  assign n707 = n579 & n620;
  assign n708 = n493 & n707;
  assign n709 = ~n584 & n708;
  assign n710 = ~pi011 & n707;
  assign n711 = n449 & n710;
  assign n712 = ~n709 & ~n711;
  assign n713 = ~n706 & n712;
  assign n714 = n292 & ~n360;
  assign n715 = n644 & n714;
  assign n716 = ~n698 & ~n715;
  assign n717 = n507 & n567;
  assign n718 = ~n716 & n717;
  assign n719 = n405 & n551;
  assign n720 = pi006 & ~n687;
  assign n721 = n719 & n720;
  assign n722 = ~n442 & ~n493;
  assign n723 = n443 & n549;
  assign n724 = ~n722 & n723;
  assign n725 = ~pi014 & n319;
  assign n726 = n687 & n725;
  assign n727 = pi006 & ~pi012;
  assign n728 = n726 & n727;
  assign n729 = ~n724 & ~n728;
  assign n730 = n349 & n519;
  assign n731 = n314 & n730;
  assign n732 = n334 & n335;
  assign n733 = n314 & n732;
  assign n734 = ~pi006 & n733;
  assign n735 = n549 & n725;
  assign n736 = n332 & n735;
  assign n737 = ~pi027 & pi028;
  assign n738 = ~pi024 & ~pi029;
  assign n739 = n327 & n738;
  assign n740 = n737 & n739;
  assign n741 = n340 & n672;
  assign n742 = n349 & n454;
  assign n743 = ~pi002 & n295;
  assign n744 = pi000 & n743;
  assign n745 = ~pi112 & n742;
  assign n746 = n744 & n745;
  assign n747 = pi001 & pi006;
  assign n748 = n518 & n747;
  assign n749 = n744 & n748;
  assign n750 = ~n746 & ~n749;
  assign n751 = n311 & n349;
  assign n752 = n376 & n751;
  assign n753 = n369 & n498;
  assign n754 = ~pi110 & n376;
  assign n755 = n753 & n754;
  assign n756 = ~pi001 & n376;
  assign n757 = n500 & n756;
  assign n758 = n335 & n498;
  assign n759 = ~pi118 & n758;
  assign n760 = n376 & n759;
  assign n761 = n493 & n725;
  assign n762 = pi015 & n761;
  assign n763 = n549 & n762;
  assign n764 = ~n755 & ~n757;
  assign n765 = ~n760 & n764;
  assign n766 = ~n763 & n765;
  assign n767 = ~n741 & ~n752;
  assign n768 = n750 & n767;
  assign n769 = n766 & n768;
  assign n770 = n740 & ~n769;
  assign n771 = ~pi029 & n328;
  assign n772 = ~pi019 & n418;
  assign n773 = ~pi016 & n772;
  assign n774 = n596 & n773;
  assign n775 = n416 & n774;
  assign n776 = ~pi016 & ~pi019;
  assign n777 = n376 & n776;
  assign n778 = n426 & n777;
  assign n779 = n596 & n778;
  assign n780 = ~n775 & ~n779;
  assign n781 = pi005 & n520;
  assign n782 = ~pi004 & n781;
  assign n783 = n780 & ~n782;
  assign n784 = n771 & ~n783;
  assign n785 = ~pi008 & ~pi014;
  assign n786 = n308 & n351;
  assign n787 = n785 & n786;
  assign n788 = n290 & n787;
  assign n789 = n303 & n493;
  assign n790 = n788 & n789;
  assign n791 = ~n360 & n492;
  assign n792 = n790 & n791;
  assign n793 = n292 & n311;
  assign n794 = n349 & n793;
  assign n795 = ~n360 & n794;
  assign n796 = ~n792 & ~n795;
  assign n797 = n479 & n520;
  assign n798 = ~pi029 & n408;
  assign n799 = ~n330 & ~n798;
  assign n800 = ~pi024 & ~pi027;
  assign n801 = n327 & n800;
  assign n802 = ~pi029 & n801;
  assign n803 = n799 & ~n802;
  assign n804 = n797 & ~n803;
  assign n805 = n796 & ~n804;
  assign n806 = ~n784 & n805;
  assign n807 = n388 & n773;
  assign n808 = pi108 & ~pi109;
  assign n809 = n487 & n566;
  assign n810 = n293 & n809;
  assign n811 = ~pi045 & ~pi122;
  assign n812 = n810 & n811;
  assign n813 = n808 & n812;
  assign n814 = n347 & n813;
  assign n815 = pi045 & n808;
  assign n816 = ~pi122 & ~n815;
  assign n817 = pi108 & n816;
  assign n818 = n347 & n810;
  assign n819 = ~n817 & n818;
  assign n820 = ~n814 & ~n819;
  assign n821 = ~n807 & n820;
  assign n822 = n492 & ~n821;
  assign n823 = pi014 & n339;
  assign n824 = n493 & n823;
  assign n825 = n405 & n492;
  assign n826 = ~n311 & ~n825;
  assign n827 = n349 & n549;
  assign n828 = ~pi108 & ~pi122;
  assign n829 = n827 & n828;
  assign n830 = ~n826 & n829;
  assign n831 = ~pi122 & ~n808;
  assign n832 = n827 & ~n831;
  assign n833 = ~pi049 & n500;
  assign n834 = ~n498 & ~n833;
  assign n835 = ~n825 & n834;
  assign n836 = n832 & ~n835;
  assign n837 = n606 & n628;
  assign n838 = ~pi043 & ~pi068;
  assign n839 = ~pi044 & ~pi067;
  assign n840 = pi042 & n838;
  assign n841 = n839 & n840;
  assign n842 = n837 & n841;
  assign n843 = ~pi042 & n837;
  assign n844 = pi044 & pi067;
  assign n845 = n838 & n844;
  assign n846 = n843 & n845;
  assign n847 = pi043 & pi068;
  assign n848 = n839 & n847;
  assign n849 = n843 & n848;
  assign n850 = ~n846 & ~n849;
  assign n851 = ~n842 & n850;
  assign n852 = n493 & n580;
  assign n853 = n290 & n457;
  assign n854 = pi014 & n853;
  assign n855 = n852 & n854;
  assign n856 = ~pi054 & ~n492;
  assign n857 = n855 & ~n856;
  assign n858 = n851 & ~n857;
  assign n859 = n465 & n682;
  assign n860 = n625 & n859;
  assign n861 = n858 & ~n860;
  assign n862 = ~pi007 & n465;
  assign n863 = n300 & n862;
  assign n864 = n585 & n863;
  assign n865 = n370 & n500;
  assign n866 = ~pi119 & n758;
  assign n867 = n335 & n500;
  assign n868 = ~n866 & ~n867;
  assign n869 = n572 & ~n868;
  assign n870 = pi029 & n869;
  assign n871 = ~n865 & ~n870;
  assign n872 = ~n864 & n871;
  assign n873 = n567 & n813;
  assign n874 = pi049 & n500;
  assign n875 = ~pi051 & n874;
  assign n876 = n832 & n875;
  assign n877 = ~n873 & ~n876;
  assign n878 = ~pi021 & n810;
  assign n879 = ~pi022 & n878;
  assign n880 = ~n817 & n879;
  assign n881 = n877 & ~n880;
  assign n882 = n872 & n881;
  assign n883 = ~pi018 & n347;
  assign n884 = ~pi020 & n353;
  assign n885 = n883 & n884;
  assign n886 = n361 & n885;
  assign n887 = ~pi017 & n886;
  assign n888 = ~n824 & ~n830;
  assign n889 = ~n836 & n888;
  assign n890 = ~n887 & n889;
  assign n891 = n806 & n890;
  assign n892 = ~n822 & n891;
  assign n893 = n861 & n882;
  assign n894 = n892 & n893;
  assign n895 = pi101 & ~pi102;
  assign n896 = pi103 & n895;
  assign n897 = n609 & n862;
  assign n898 = n493 & n584;
  assign n899 = n897 & n898;
  assign n900 = ~pi007 & n675;
  assign n901 = n609 & n900;
  assign n902 = pi012 & n303;
  assign n903 = n901 & n902;
  assign n904 = pi013 & n903;
  assign n905 = ~n899 & ~n904;
  assign n906 = n896 & ~n905;
  assign n907 = n798 & n906;
  assign n908 = ~n721 & ~n731;
  assign n909 = ~n734 & n908;
  assign n910 = ~n736 & n909;
  assign n911 = n729 & n910;
  assign n912 = ~n629 & n663;
  assign n913 = ~n666 & n912;
  assign n914 = ~n574 & n911;
  assign n915 = ~n624 & n651;
  assign n916 = ~n671 & n915;
  assign n917 = n913 & n914;
  assign n918 = n701 & n713;
  assign n919 = ~n718 & n918;
  assign n920 = n916 & n917;
  assign n921 = n696 & ~n770;
  assign n922 = n920 & n921;
  assign n923 = n619 & n919;
  assign n924 = ~n907 & n923;
  assign n925 = n922 & n924;
  assign n926 = n565 & n925;
  assign po000 = ~n894 | ~n926;
  assign n928 = pi022 & n361;
  assign n929 = ~pi021 & n928;
  assign n930 = pi018 & n599;
  assign n931 = ~pi020 & n930;
  assign n932 = n929 & n931;
  assign n933 = ~pi018 & n567;
  assign n934 = n390 & n933;
  assign n935 = n361 & n934;
  assign n936 = ~pi019 & n935;
  assign n937 = n644 & n717;
  assign n938 = ~n360 & n416;
  assign n939 = n937 & n938;
  assign n940 = ~n936 & ~n939;
  assign n941 = n619 & n940;
  assign n942 = n740 & n906;
  assign n943 = ~pi007 & n607;
  assign n944 = n300 & n943;
  assign n945 = n581 & n944;
  assign n946 = ~n942 & ~n945;
  assign n947 = n623 & ~n678;
  assign n948 = n442 & ~n947;
  assign n949 = n419 & n566;
  assign n950 = n938 & n949;
  assign n951 = n510 & n950;
  assign n952 = pi019 & n951;
  assign n953 = ~pi023 & n952;
  assign n954 = n375 & n529;
  assign n955 = ~pi002 & n954;
  assign n956 = n518 & n955;
  assign n957 = pi005 & pi006;
  assign n958 = n719 & n957;
  assign n959 = pi007 & n465;
  assign n960 = ~pi014 & n437;
  assign n961 = n959 & n960;
  assign n962 = n330 & n961;
  assign n963 = n332 & n580;
  assign n964 = n962 & n963;
  assign n965 = ~pi015 & n332;
  assign n966 = n314 & n725;
  assign n967 = ~pi006 & n965;
  assign n968 = n966 & n967;
  assign n969 = n809 & n928;
  assign n970 = pi001 & pi003;
  assign n971 = n310 & n970;
  assign n972 = ~pi021 & n566;
  assign n973 = ~pi019 & ~pi023;
  assign n974 = n419 & n973;
  assign n975 = n972 & n974;
  assign n976 = ~n971 & ~n975;
  assign n977 = n938 & ~n976;
  assign n978 = ~n956 & ~n958;
  assign n979 = ~n968 & n978;
  assign n980 = ~n684 & n979;
  assign n981 = ~n670 & ~n969;
  assign n982 = n980 & n981;
  assign n983 = ~n932 & ~n964;
  assign n984 = ~n977 & n983;
  assign n985 = ~n948 & n982;
  assign n986 = ~n953 & n985;
  assign n987 = n984 & n986;
  assign n988 = n941 & n987;
  assign n989 = n946 & n988;
  assign n990 = ~n330 & ~n740;
  assign n991 = ~n741 & ~n763;
  assign n992 = ~pi122 & n349;
  assign n993 = n376 & n992;
  assign n994 = ~pi108 & n993;
  assign n995 = n311 & n994;
  assign n996 = n991 & ~n995;
  assign n997 = pi122 & n752;
  assign n998 = ~pi007 & n757;
  assign n999 = ~n759 & ~n867;
  assign n1000 = n307 & ~n999;
  assign n1001 = ~n755 & ~n998;
  assign n1002 = ~n1000 & n1001;
  assign n1003 = n996 & ~n997;
  assign n1004 = n1002 & n1003;
  assign n1005 = ~n990 & ~n1004;
  assign n1006 = ~pi013 & ~pi014;
  assign n1007 = ~pi012 & ~pi015;
  assign n1008 = n677 & n1007;
  assign n1009 = ~n1006 & n1008;
  assign n1010 = n663 & ~n1009;
  assign n1011 = n449 & n703;
  assign n1012 = pi008 & n1011;
  assign n1013 = ~n789 & ~n1012;
  assign n1014 = n859 & ~n1013;
  assign n1015 = n606 & n665;
  assign n1016 = n302 & n726;
  assign n1017 = pi015 & n1016;
  assign n1018 = ~pi006 & n1017;
  assign n1019 = pi108 & n307;
  assign n1020 = n751 & ~n990;
  assign n1021 = n1019 & n1020;
  assign n1022 = ~n1015 & ~n1021;
  assign n1023 = ~n1018 & n1022;
  assign n1024 = ~pi013 & n628;
  assign n1025 = ~pi011 & n1024;
  assign n1026 = pi013 & n728;
  assign n1027 = pi020 & n482;
  assign n1028 = n930 & n1027;
  assign n1029 = n416 & n1028;
  assign n1030 = pi029 & n537;
  assign n1031 = n1029 & n1030;
  assign n1032 = pi013 & n723;
  assign n1033 = ~pi015 & n302;
  assign n1034 = ~n332 & ~n1033;
  assign n1035 = n735 & ~n1034;
  assign n1036 = n417 & n642;
  assign n1037 = ~n643 & ~n1036;
  assign n1038 = n778 & ~n1037;
  assign n1039 = ~n689 & ~n734;
  assign n1040 = ~n1032 & ~n1035;
  assign n1041 = ~n1038 & n1040;
  assign n1042 = n1039 & n1041;
  assign n1043 = ~n1031 & n1042;
  assign n1044 = n672 & n678;
  assign n1045 = n442 & n665;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = n361 & n630;
  assign n1048 = n974 & n1047;
  assign n1049 = n390 & n485;
  assign n1050 = n516 & n1049;
  assign n1051 = ~n1048 & ~n1050;
  assign n1052 = n330 & ~n750;
  assign n1053 = ~pi108 & n308;
  assign n1054 = pi109 & n1053;
  assign n1055 = n330 & n1054;
  assign n1056 = n740 & n1053;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = n751 & ~n1057;
  assign n1059 = ~n307 & n556;
  assign n1060 = n401 & n596;
  assign n1061 = n361 & n1060;
  assign n1062 = ~pi019 & n1061;
  assign n1063 = ~n631 & ~n1062;
  assign n1064 = ~pi022 & n359;
  assign n1065 = pi019 & n390;
  assign n1066 = n361 & n1065;
  assign n1067 = n1064 & n1066;
  assign n1068 = n1063 & ~n1067;
  assign n1069 = pi018 & ~pi021;
  assign n1070 = pi020 & pi022;
  assign n1071 = n1069 & n1070;
  assign n1072 = n698 & n1071;
  assign n1073 = n351 & n636;
  assign n1074 = n638 & n642;
  assign n1075 = n1073 & n1074;
  assign n1076 = ~pi022 & n507;
  assign n1077 = n974 & n1076;
  assign n1078 = ~n1075 & ~n1077;
  assign n1079 = n361 & ~n1078;
  assign n1080 = pi017 & n352;
  assign n1081 = n566 & n1080;
  assign n1082 = n482 & n598;
  assign n1083 = n361 & n1082;
  assign n1084 = n1081 & n1083;
  assign n1085 = ~pi025 & n738;
  assign n1086 = n737 & n1085;
  assign n1087 = n1029 & n1086;
  assign n1088 = pi026 & n1087;
  assign n1089 = n314 & n493;
  assign n1090 = n725 & n1089;
  assign n1091 = ~pi006 & n1090;
  assign n1092 = n416 & ~n571;
  assign n1093 = pi029 & n328;
  assign n1094 = pi027 & pi028;
  assign n1095 = n739 & n1094;
  assign n1096 = ~n1093 & ~n1095;
  assign n1097 = n1092 & ~n1096;
  assign n1098 = ~n1084 & ~n1091;
  assign n1099 = ~n1097 & n1098;
  assign n1100 = ~n1088 & n1099;
  assign n1101 = n894 & n1100;
  assign n1102 = n507 & n974;
  assign n1103 = n483 & n1102;
  assign n1104 = ~n360 & n1103;
  assign n1105 = ~n641 & ~n1059;
  assign n1106 = ~n432 & n1105;
  assign n1107 = ~n1014 & ~n1026;
  assign n1108 = ~n1052 & ~n1058;
  assign n1109 = n1107 & n1108;
  assign n1110 = n1051 & n1106;
  assign n1111 = n1109 & n1110;
  assign n1112 = ~n423 & n1010;
  assign n1113 = ~n1025 & n1046;
  assign n1114 = ~n1072 & ~n1079;
  assign n1115 = ~n1104 & n1114;
  assign n1116 = n1112 & n1113;
  assign n1117 = n1023 & n1111;
  assign n1118 = n1068 & n1117;
  assign n1119 = n1115 & n1116;
  assign n1120 = n1043 & n1119;
  assign n1121 = ~n1005 & n1118;
  assign n1122 = n1120 & n1121;
  assign n1123 = n548 & n1122;
  assign n1124 = n989 & n1123;
  assign po001 = ~n1101 | ~n1124;
  assign n1126 = n302 & n373;
  assign po002 = ~pi015 & n1126;
  assign n1128 = n315 & n349;
  assign n1129 = n744 & n1128;
  assign n1130 = ~pi115 & n1129;
  assign n1131 = pi112 & ~pi123;
  assign n1132 = n1130 & n1131;
  assign n1133 = n492 & n1132;
  assign n1134 = ~pi056 & pi122;
  assign n1135 = pi055 & n1134;
  assign n1136 = ~pi044 & pi055;
  assign n1137 = n345 & ~n1136;
  assign n1138 = ~n1135 & ~n1137;
  assign n1139 = pi035 & ~pi123;
  assign n1140 = ~pi112 & n1130;
  assign n1141 = n306 & n744;
  assign n1142 = ~pi112 & n1141;
  assign n1143 = n314 & n1142;
  assign n1144 = ~n1140 & ~n1143;
  assign n1145 = ~n1139 & ~n1144;
  assign n1146 = ~pi079 & ~pi123;
  assign n1147 = ~pi046 & n1142;
  assign n1148 = n293 & n1147;
  assign n1149 = ~pi031 & n1146;
  assign n1150 = n1148 & n1149;
  assign n1151 = ~n1145 & ~n1150;
  assign n1152 = n687 & n744;
  assign n1153 = n349 & n1152;
  assign n1154 = n1151 & ~n1153;
  assign n1155 = ~n1138 & ~n1154;
  assign n1156 = ~n1133 & ~n1155;
  assign n1157 = ~pi079 & n1148;
  assign n1158 = pi122 & n1138;
  assign n1159 = pi123 & ~n1158;
  assign n1160 = n1157 & n1159;
  assign n1161 = n376 & n933;
  assign n1162 = pi020 & n1161;
  assign n1163 = n390 & n973;
  assign n1164 = n1162 & n1163;
  assign n1165 = n345 & n1164;
  assign n1166 = n992 & n1152;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~pi031 & ~pi122;
  assign n1169 = n1157 & n1168;
  assign n1170 = pi003 & n349;
  assign n1171 = n316 & n1170;
  assign n1172 = pi002 & n1171;
  assign n1173 = pi065 & ~pi112;
  assign n1174 = n293 & n1173;
  assign n1175 = n1172 & n1174;
  assign n1176 = ~pi122 & n1175;
  assign n1177 = n333 & n475;
  assign n1178 = pi061 & n1177;
  assign n1179 = n296 & n992;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = pi112 & n293;
  assign n1182 = ~n1180 & n1181;
  assign n1183 = ~n1176 & ~n1182;
  assign n1184 = ~n1169 & n1183;
  assign n1185 = ~n549 & ~n1174;
  assign n1186 = n1172 & ~n1185;
  assign n1187 = ~n1138 & n1186;
  assign n1188 = pi001 & n296;
  assign n1189 = pi061 & n1188;
  assign n1190 = ~pi061 & pi065;
  assign n1191 = n1177 & n1190;
  assign n1192 = ~n1189 & ~n1191;
  assign n1193 = ~pi112 & ~n1192;
  assign n1194 = n293 & n1193;
  assign n1195 = ~n1158 & n1194;
  assign n1196 = n549 & n1179;
  assign n1197 = ~n1187 & ~n1196;
  assign n1198 = ~n1195 & n1197;
  assign n1199 = ~pi122 & n1145;
  assign n1200 = n292 & n425;
  assign n1201 = n376 & n1141;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1158 & ~n1202;
  assign n1204 = ~pi035 & pi112;
  assign n1205 = ~pi123 & n1204;
  assign n1206 = n314 & n1205;
  assign n1207 = n1141 & n1206;
  assign n1208 = ~n1203 & ~n1207;
  assign n1209 = ~n1199 & n1208;
  assign n1210 = ~n1160 & n1167;
  assign n1211 = n1198 & n1210;
  assign n1212 = n1184 & n1209;
  assign n1213 = n1211 & n1212;
  assign po003 = ~n1156 | ~n1213;
  assign n1215 = n746 & n798;
  assign n1216 = ~n1138 & n1215;
  assign n1217 = ~pi008 & n579;
  assign n1218 = n786 & n1217;
  assign n1219 = n702 & n1218;
  assign n1220 = ~n749 & ~n1219;
  assign n1221 = n798 & ~n1220;
  assign n1222 = ~n1158 & n1221;
  assign n1223 = ~n1216 & ~n1222;
  assign n1224 = n304 & n1218;
  assign n1225 = ~pi047 & n1224;
  assign n1226 = pi122 & n1225;
  assign n1227 = n330 & n1226;
  assign n1228 = pi027 & n1093;
  assign n1229 = ~n746 & n1220;
  assign n1230 = n1228 & ~n1229;
  assign n1231 = ~pi122 & n1215;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1227 & n1232;
  assign n1234 = n492 & ~n1138;
  assign n1235 = n1225 & n1234;
  assign n1236 = n1233 & ~n1235;
  assign n1237 = pi079 & ~n1158;
  assign n1238 = n1148 & n1237;
  assign n1239 = n1223 & ~n1238;
  assign po004 = ~n1236 | ~n1239;
  assign n1241 = pi022 & n315;
  assign n1242 = n417 & n1241;
  assign n1243 = n362 & n973;
  assign n1244 = ~n360 & n1243;
  assign n1245 = n1242 & n1244;
  assign n1246 = n376 & n974;
  assign n1247 = n630 & n1246;
  assign n1248 = n315 & n1028;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = ~n801 & ~n1249;
  assign n1251 = ~po002 & ~n1250;
  assign n1252 = ~pi027 & ~pi028;
  assign n1253 = ~pi026 & n1252;
  assign n1254 = ~pi007 & n960;
  assign n1255 = n465 & n1254;
  assign n1256 = ~n1253 & n1255;
  assign n1257 = n450 & n1256;
  assign n1258 = ~pi022 & n566;
  assign n1259 = n592 & n1258;
  assign n1260 = pi021 & pi023;
  assign n1261 = n1259 & n1260;
  assign n1262 = n416 & n1261;
  assign n1263 = pi028 & ~pi029;
  assign n1264 = ~n801 & n1263;
  assign n1265 = n1262 & n1264;
  assign n1266 = ~n1257 & ~n1265;
  assign n1267 = n798 & n1172;
  assign n1268 = n416 & n1267;
  assign n1269 = ~n360 & n1268;
  assign n1270 = n518 & n798;
  assign n1271 = n1177 & n1270;
  assign n1272 = ~n360 & n1271;
  assign n1273 = ~n1269 & ~n1272;
  assign n1274 = pi061 & ~n1273;
  assign n1275 = n362 & n485;
  assign n1276 = n315 & n482;
  assign n1277 = n1275 & n1276;
  assign n1278 = n667 & n1277;
  assign n1279 = ~n344 & n1278;
  assign n1280 = n351 & n453;
  assign n1281 = ~n1158 & n1280;
  assign n1282 = n416 & ~n1253;
  assign n1283 = n1243 & n1282;
  assign n1284 = pi021 & n566;
  assign n1285 = n1283 & n1284;
  assign n1286 = ~pi022 & n1285;
  assign n1287 = ~n1245 & ~n1281;
  assign n1288 = ~n1274 & n1287;
  assign n1289 = ~n1279 & ~n1286;
  assign n1290 = n1288 & n1289;
  assign n1291 = n1266 & n1290;
  assign po008 = ~n1251 | ~n1291;
  assign n1293 = ~pi061 & ~n1273;
  assign n1294 = n376 & n1188;
  assign n1295 = n389 & n667;
  assign n1296 = pi023 & n637;
  assign n1297 = n1295 & n1296;
  assign n1298 = ~pi035 & n1297;
  assign n1299 = ~pi036 & n1298;
  assign n1300 = n567 & n1299;
  assign n1301 = ~pi037 & n1300;
  assign n1302 = ~n360 & n1301;
  assign n1303 = ~n1294 & ~n1302;
  assign n1304 = pi027 & n535;
  assign n1305 = pi029 & n1304;
  assign n1306 = pi026 & n1305;
  assign n1307 = ~n1303 & n1306;
  assign n1308 = n1085 & n1094;
  assign n1309 = pi061 & n1294;
  assign n1310 = pi026 & n1309;
  assign n1311 = n1308 & n1310;
  assign n1312 = ~n1307 & ~n1311;
  assign n1313 = pi037 & n1299;
  assign n1314 = n347 & n1313;
  assign n1315 = ~n1300 & ~n1314;
  assign n1316 = ~n360 & ~n1315;
  assign n1317 = ~n740 & ~n1228;
  assign n1318 = ~n1030 & n1317;
  assign n1319 = n1316 & ~n1318;
  assign n1320 = n1312 & ~n1319;
  assign n1321 = n798 & n1092;
  assign n1322 = n573 & ~n602;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = n1320 & n1323;
  assign n1325 = n303 & n332;
  assign n1326 = n1255 & n1325;
  assign n1327 = pi029 & n1326;
  assign n1328 = n515 & n1163;
  assign n1329 = ~n990 & n1328;
  assign n1330 = pi031 & ~pi079;
  assign n1331 = ~pi123 & n1330;
  assign n1332 = ~pi035 & n1331;
  assign n1333 = n1148 & n1332;
  assign n1334 = n798 & n1333;
  assign n1335 = n896 & n903;
  assign n1336 = ~pi013 & n1335;
  assign n1337 = n491 & n535;
  assign n1338 = pi026 & n1337;
  assign n1339 = n1336 & n1338;
  assign n1340 = ~n1334 & ~n1339;
  assign n1341 = ~n1329 & n1340;
  assign n1342 = ~pi035 & pi036;
  assign n1343 = ~pi022 & n637;
  assign n1344 = n1295 & n1343;
  assign n1345 = n1342 & n1344;
  assign n1346 = pi023 & n360;
  assign n1347 = ~n1317 & ~n1346;
  assign n1348 = n1345 & n1347;
  assign n1349 = n1341 & ~n1348;
  assign n1350 = ~n1327 & n1349;
  assign n1351 = n480 & n601;
  assign n1352 = n593 & n667;
  assign n1353 = n347 & n1352;
  assign n1354 = ~n1351 & ~n1353;
  assign n1355 = ~pi039 & ~n360;
  assign n1356 = ~n1354 & n1355;
  assign n1357 = n480 & n798;
  assign n1358 = ~n687 & ~n1357;
  assign n1359 = n955 & ~n1358;
  assign n1360 = n938 & n972;
  assign n1361 = n575 & n928;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = n507 & n928;
  assign n1364 = n1362 & ~n1363;
  assign n1365 = ~pi019 & pi023;
  assign n1366 = n419 & n1365;
  assign n1367 = ~n1364 & n1366;
  assign n1368 = ~n360 & n788;
  assign n1369 = ~n302 & n580;
  assign n1370 = n1368 & n1369;
  assign n1371 = n347 & n566;
  assign n1372 = ~pi019 & n1371;
  assign n1373 = n363 & n1372;
  assign n1374 = ~n1370 & ~n1373;
  assign n1375 = n329 & ~n360;
  assign n1376 = pi029 & n1375;
  assign n1377 = ~n740 & ~n1376;
  assign n1378 = ~pi021 & n315;
  assign n1379 = n434 & n1378;
  assign n1380 = pi019 & n362;
  assign n1381 = n1379 & n1380;
  assign n1382 = ~n1377 & n1381;
  assign n1383 = pi023 & n952;
  assign n1384 = n773 & n1284;
  assign n1385 = ~n360 & n376;
  assign n1386 = n1384 & n1385;
  assign n1387 = ~pi023 & n354;
  assign n1388 = n972 & n1387;
  assign n1389 = n361 & n1388;
  assign n1390 = ~n1386 & ~n1389;
  assign n1391 = pi022 & ~n1390;
  assign n1392 = pi020 & n599;
  assign n1393 = n483 & n1392;
  assign n1394 = pi018 & n1393;
  assign n1395 = ~n360 & n1394;
  assign n1396 = pi002 & n309;
  assign n1397 = ~pi003 & n1396;
  assign n1398 = ~n404 & ~n1397;
  assign n1399 = pi001 & ~n360;
  assign n1400 = ~pi006 & ~pi007;
  assign n1401 = n687 & n1400;
  assign n1402 = n1399 & n1401;
  assign n1403 = ~n1398 & n1402;
  assign n1404 = n361 & n567;
  assign n1405 = ~pi020 & n1387;
  assign n1406 = n1404 & n1405;
  assign n1407 = ~n1403 & ~n1406;
  assign n1408 = ~n1383 & n1407;
  assign n1409 = ~n1395 & n1408;
  assign n1410 = ~n1391 & n1409;
  assign n1411 = ~n1367 & ~n1382;
  assign n1412 = n1374 & n1411;
  assign n1413 = n1410 & n1412;
  assign n1414 = ~n1356 & ~n1359;
  assign n1415 = n1413 & n1414;
  assign n1416 = n308 & n444;
  assign n1417 = ~n302 & n1416;
  assign n1418 = n362 & n667;
  assign n1419 = pi023 & n1418;
  assign n1420 = n483 & n1419;
  assign n1421 = ~n360 & n1420;
  assign n1422 = ~n1417 & ~n1421;
  assign n1423 = ~n668 & ~n1284;
  assign n1424 = n419 & ~n1423;
  assign n1425 = n667 & n1080;
  assign n1426 = pi022 & n1425;
  assign n1427 = ~n1424 & ~n1426;
  assign n1428 = ~pi023 & n938;
  assign n1429 = ~n1427 & n1428;
  assign n1430 = n1422 & ~n1429;
  assign n1431 = n338 & n744;
  assign n1432 = ~n360 & n1431;
  assign n1433 = n1430 & ~n1432;
  assign n1434 = pi047 & pi113;
  assign n1435 = n1224 & n1434;
  assign n1436 = n345 & n1435;
  assign n1437 = ~pi061 & ~pi065;
  assign n1438 = ~pi112 & n1437;
  assign n1439 = n293 & n1438;
  assign n1440 = n1188 & n1439;
  assign n1441 = ~n474 & n1440;
  assign n1442 = ~n1436 & ~n1441;
  assign n1443 = n330 & ~n1442;
  assign n1444 = n334 & n756;
  assign n1445 = ~n360 & n1444;
  assign n1446 = ~n899 & ~n903;
  assign n1447 = pi029 & ~n1252;
  assign n1448 = n327 & ~n1447;
  assign n1449 = n360 & ~n1448;
  assign n1450 = n896 & ~n1449;
  assign n1451 = ~n1446 & ~n1450;
  assign n1452 = n360 & n1094;
  assign n1453 = ~n905 & n1452;
  assign n1454 = ~n1451 & ~n1453;
  assign n1455 = pi122 & n740;
  assign n1456 = n1435 & n1455;
  assign n1457 = ~n1445 & ~n1456;
  assign n1458 = n1454 & n1457;
  assign n1459 = ~n1443 & n1458;
  assign n1460 = n1433 & n1459;
  assign n1461 = pi046 & n1141;
  assign n1462 = n293 & n1461;
  assign n1463 = pi035 & n1344;
  assign n1464 = n585 & n897;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~pi079 & n1139;
  assign n1467 = ~n1332 & ~n1466;
  assign n1468 = n1148 & ~n1467;
  assign n1469 = n1465 & ~n1468;
  assign n1470 = ~n1462 & n1469;
  assign n1471 = n1376 & ~n1470;
  assign n1472 = n896 & ~n1446;
  assign n1473 = ~n360 & n1228;
  assign n1474 = n1472 & n1473;
  assign n1475 = n511 & n1049;
  assign n1476 = n317 & n452;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = n416 & ~n1477;
  assign n1479 = n438 & n862;
  assign n1480 = n304 & n1479;
  assign n1481 = ~n1478 & ~n1480;
  assign n1482 = n315 & n601;
  assign n1483 = n1481 & ~n1482;
  assign n1484 = n1264 & ~n1483;
  assign n1485 = ~pi001 & n744;
  assign n1486 = n314 & ~n360;
  assign n1487 = ~pi007 & n1486;
  assign n1488 = ~n361 & ~n1487;
  assign n1489 = n1485 & ~n1488;
  assign n1490 = n386 & n487;
  assign n1491 = n596 & n1387;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = n938 & ~n1492;
  assign n1494 = n384 & n938;
  assign n1495 = n1405 & n1494;
  assign n1496 = ~n1489 & ~n1495;
  assign n1497 = ~n1493 & n1496;
  assign n1498 = ~n1095 & ~n1338;
  assign n1499 = n1029 & ~n1498;
  assign n1500 = n483 & n1243;
  assign n1501 = n667 & n1500;
  assign n1502 = n537 & n1501;
  assign n1503 = ~n1499 & ~n1502;
  assign n1504 = n798 & n1500;
  assign n1505 = n566 & n1504;
  assign n1506 = n592 & n1379;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n360 & ~n1507;
  assign n1509 = n1503 & ~n1508;
  assign n1510 = n1401 & n1485;
  assign n1511 = ~n1253 & n1510;
  assign n1512 = pi029 & ~pi061;
  assign n1513 = n549 & n1177;
  assign n1514 = n537 & ~n1512;
  assign n1515 = n1513 & n1514;
  assign n1516 = n315 & n592;
  assign n1517 = ~pi045 & n740;
  assign n1518 = ~n1376 & ~n1517;
  assign n1519 = n630 & ~n1518;
  assign n1520 = n1516 & n1519;
  assign n1521 = n1139 & ~n1144;
  assign n1522 = ~n1518 & n1521;
  assign n1523 = pi022 & n1284;
  assign n1524 = n1283 & n1523;
  assign n1525 = pi015 & n302;
  assign n1526 = n373 & n1525;
  assign n1527 = pi023 & n482;
  assign n1528 = n950 & n1527;
  assign n1529 = pi045 & ~pi056;
  assign n1530 = pi115 & n1129;
  assign n1531 = ~pi044 & pi045;
  assign n1532 = pi056 & ~n1531;
  assign n1533 = ~n1529 & ~n1532;
  assign n1534 = n329 & n1533;
  assign n1535 = n1530 & n1534;
  assign n1536 = ~pi029 & n1535;
  assign n1537 = ~n1528 & ~n1536;
  assign n1538 = n304 & n1256;
  assign n1539 = ~pi023 & n1065;
  assign n1540 = n717 & n1539;
  assign n1541 = n1282 & n1540;
  assign n1542 = ~n1511 & ~n1515;
  assign n1543 = ~n1526 & n1542;
  assign n1544 = ~n1520 & n1543;
  assign n1545 = ~n1524 & n1544;
  assign n1546 = ~n1293 & ~n1522;
  assign n1547 = n1537 & ~n1541;
  assign n1548 = n1546 & n1547;
  assign n1549 = ~n1538 & n1545;
  assign n1550 = n1548 & n1549;
  assign n1551 = ~n1474 & n1497;
  assign n1552 = n1550 & n1551;
  assign n1553 = ~n1471 & ~n1484;
  assign n1554 = n1509 & n1553;
  assign n1555 = n1552 & n1554;
  assign n1556 = n1350 & n1555;
  assign n1557 = n1415 & n1460;
  assign n1558 = n1556 & n1557;
  assign po009 = ~n1324 | ~n1558;
  assign n1560 = pi020 & n935;
  assign n1561 = pi007 & n500;
  assign n1562 = n349 & n498;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = ~n759 & n1563;
  assign n1565 = ~pi109 & n1056;
  assign n1566 = ~n1564 & n1565;
  assign n1567 = pi027 & n739;
  assign n1568 = pi025 & pi056;
  assign n1569 = n344 & n1568;
  assign n1570 = ~n1567 & ~n1569;
  assign n1571 = n403 & n744;
  assign n1572 = ~n1570 & n1571;
  assign n1573 = ~n1038 & ~n1572;
  assign n1574 = ~n1566 & n1573;
  assign n1575 = n1323 & n1574;
  assign n1576 = n334 & n337;
  assign n1577 = n322 & n1576;
  assign n1578 = ~pi005 & n1577;
  assign n1579 = n426 & n1296;
  assign n1580 = n596 & n1579;
  assign n1581 = pi072 & n1580;
  assign n1582 = n426 & n637;
  assign n1583 = n1036 & n1582;
  assign n1584 = n740 & n1583;
  assign n1585 = ~pi031 & ~pi034;
  assign n1586 = n315 & n498;
  assign n1587 = pi007 & n1585;
  assign n1588 = n1586 & n1587;
  assign n1589 = ~n1584 & ~n1588;
  assign n1590 = n418 & n636;
  assign n1591 = n1360 & n1590;
  assign n1592 = n304 & n678;
  assign n1593 = ~n1338 & ~n1567;
  assign n1594 = n1029 & ~n1593;
  assign n1595 = n340 & n494;
  assign n1596 = n494 & n735;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = n310 & n315;
  assign n1599 = n350 & n1598;
  assign n1600 = pi039 & n1599;
  assign n1601 = n1597 & ~n1600;
  assign n1602 = n1585 & ~n1601;
  assign n1603 = ~n677 & ~n944;
  assign n1604 = n581 & ~n1603;
  assign n1605 = ~n1578 & ~n1591;
  assign n1606 = ~n1052 & n1605;
  assign n1607 = ~n1581 & ~n1592;
  assign n1608 = n1606 & n1607;
  assign n1609 = ~n1045 & ~n1560;
  assign n1610 = n1589 & n1609;
  assign n1611 = ~n952 & n1608;
  assign n1612 = ~n1602 & ~n1604;
  assign n1613 = n1611 & n1612;
  assign n1614 = ~n1594 & n1610;
  assign n1615 = n1613 & n1614;
  assign po011 = ~n1575 | ~n1615;
  assign n1617 = ~n783 & n1228;
  assign n1618 = ~pi054 & n855;
  assign n1619 = n330 & n1618;
  assign n1620 = n315 & n330;
  assign n1621 = n753 & n1620;
  assign n1622 = ~n1619 & ~n1621;
  assign n1623 = n1371 & n1582;
  assign n1624 = pi021 & n667;
  assign n1625 = ~n1523 & ~n1624;
  assign n1626 = n577 & ~n1625;
  assign n1627 = ~n1623 & ~n1626;
  assign n1628 = n519 & n827;
  assign n1629 = n1627 & ~n1628;
  assign n1630 = ~n496 & n1629;
  assign n1631 = n330 & ~n1630;
  assign n1632 = n807 & n1376;
  assign n1633 = n955 & n1620;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = ~n1617 & n1634;
  assign n1636 = n1622 & ~n1631;
  assign po013 = ~n1635 | ~n1636;
  assign n1638 = ~pi023 & n1582;
  assign n1639 = n596 & n1638;
  assign n1640 = n442 & n1576;
  assign n1641 = ~n321 & n1640;
  assign n1642 = ~pi005 & n1641;
  assign n1643 = pi026 & ~n534;
  assign n1644 = n1086 & n1643;
  assign n1645 = ~n1642 & ~n1644;
  assign n1646 = ~pi090 & n1579;
  assign n1647 = ~pi091 & n1646;
  assign n1648 = ~pi092 & n1647;
  assign n1649 = n386 & n1648;
  assign n1650 = ~pi093 & n1649;
  assign n1651 = pi094 & n1650;
  assign n1652 = n789 & n1255;
  assign n1653 = n1305 & n1652;
  assign n1654 = ~pi026 & n1653;
  assign n1655 = ~n1526 & n1645;
  assign n1656 = ~n1651 & n1655;
  assign po021 = n1654 | ~n1656;
  assign po015 = n1639 | po021;
  assign n1659 = pi007 & n607;
  assign n1660 = n438 & n1659;
  assign n1661 = n580 & n1660;
  assign n1662 = n303 & n959;
  assign n1663 = n438 & n1662;
  assign n1664 = ~n1661 & ~n1663;
  assign n1665 = pi012 & ~n1664;
  assign n1666 = n492 & n1665;
  assign n1667 = n330 & n1525;
  assign n1668 = pi011 & n1667;
  assign n1669 = pi007 & pi009;
  assign n1670 = pi010 & n1669;
  assign n1671 = n960 & n1670;
  assign n1672 = n1668 & n1671;
  assign n1673 = n330 & n960;
  assign n1674 = ~pi011 & ~pi012;
  assign n1675 = n1659 & n1674;
  assign n1676 = n1673 & n1675;
  assign n1677 = pi017 & pi023;
  assign n1678 = n1073 & ~n1677;
  assign n1679 = n1242 & n1678;
  assign n1680 = ~n482 & n507;
  assign n1681 = ~pi020 & pi022;
  assign n1682 = n1069 & n1681;
  assign n1683 = ~n1680 & ~n1682;
  assign n1684 = pi016 & n315;
  assign n1685 = n772 & n1684;
  assign n1686 = ~n1683 & n1685;
  assign n1687 = n385 & n1241;
  assign n1688 = n315 & n1371;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = n1366 & ~n1689;
  assign n1691 = ~n1679 & ~n1686;
  assign n1692 = ~n1690 & n1691;
  assign n1693 = n329 & n854;
  assign n1694 = pi029 & n1693;
  assign n1695 = n304 & n1694;
  assign n1696 = pi014 & n298;
  assign n1697 = ~pi010 & n1669;
  assign n1698 = n1696 & n1697;
  assign n1699 = n438 & n1670;
  assign n1700 = n408 & n1699;
  assign n1701 = ~n1698 & ~n1700;
  assign n1702 = n332 & n653;
  assign n1703 = ~n1701 & n1702;
  assign n1704 = n437 & n1697;
  assign n1705 = pi011 & n1704;
  assign n1706 = n965 & n1705;
  assign n1707 = pi014 & n1706;
  assign n1708 = ~pi018 & pi021;
  assign n1709 = n592 & n1708;
  assign n1710 = n1385 & n1709;
  assign n1711 = n362 & n427;
  assign n1712 = ~n360 & n1711;
  assign n1713 = n883 & n1712;
  assign n1714 = ~n1710 & ~n1713;
  assign n1715 = pi023 & n315;
  assign n1716 = n1071 & n1715;
  assign n1717 = n1590 & n1716;
  assign n1718 = pi011 & n442;
  assign n1719 = n1704 & n1718;
  assign n1720 = n654 & n1671;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = n362 & n575;
  assign n1723 = n1385 & n1722;
  assign n1724 = n442 & n653;
  assign n1725 = ~pi009 & n1724;
  assign n1726 = n1254 & n1725;
  assign n1727 = n852 & n961;
  assign n1728 = pi011 & pi012;
  assign n1729 = ~pi013 & ~pi015;
  assign n1730 = n1728 & n1729;
  assign n1731 = n1254 & n1730;
  assign n1732 = n607 & n1731;
  assign n1733 = ~n1726 & ~n1727;
  assign n1734 = ~n1732 & n1733;
  assign n1735 = ~pi094 & n1650;
  assign n1736 = ~pi095 & n1735;
  assign n1737 = pi096 & n1736;
  assign n1738 = n1255 & n1702;
  assign n1739 = n330 & n1738;
  assign n1740 = n1734 & ~n1739;
  assign po020 = n1737 | ~n1740;
  assign n1742 = ~pi012 & n580;
  assign n1743 = ~n672 & ~n1742;
  assign n1744 = ~pi008 & n1698;
  assign n1745 = ~n1743 & n1744;
  assign n1746 = ~pi013 & pi015;
  assign n1747 = pi014 & ~n1746;
  assign n1748 = ~n442 & ~n1747;
  assign n1749 = n299 & n959;
  assign n1750 = ~n1748 & n1749;
  assign n1751 = n669 & n1685;
  assign n1752 = pi011 & n493;
  assign n1753 = n329 & n1699;
  assign n1754 = pi029 & n1753;
  assign n1755 = n1752 & n1754;
  assign n1756 = pi015 & n1755;
  assign n1757 = n1379 & n1590;
  assign n1758 = n652 & n962;
  assign n1759 = n299 & n1697;
  assign n1760 = n692 & n1759;
  assign n1761 = ~n1757 & ~n1760;
  assign n1762 = ~n1758 & n1761;
  assign n1763 = n362 & n1385;
  assign n1764 = n485 & n1763;
  assign n1765 = n482 & n1764;
  assign n1766 = n1027 & n1763;
  assign n1767 = n598 & n1766;
  assign n1768 = ~n1765 & ~n1767;
  assign n1769 = ~pi018 & ~n1768;
  assign n1770 = n609 & n1697;
  assign n1771 = ~pi011 & n1770;
  assign n1772 = n609 & n959;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = pi013 & ~n1773;
  assign n1775 = ~pi011 & ~pi013;
  assign n1776 = pi015 & n1775;
  assign n1777 = ~n853 & ~n1671;
  assign n1778 = n492 & n1776;
  assign n1779 = ~n1777 & n1778;
  assign n1780 = pi007 & ~pi009;
  assign n1781 = ~pi010 & ~pi011;
  assign n1782 = pi010 & pi011;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = n1780 & n1783;
  assign n1785 = pi012 & n1784;
  assign n1786 = n329 & n960;
  assign n1787 = ~pi029 & n1786;
  assign n1788 = n1785 & n1787;
  assign n1789 = n492 & n854;
  assign n1790 = ~pi013 & n1789;
  assign n1791 = ~n1671 & ~n1790;
  assign n1792 = n580 & ~n1791;
  assign n1793 = ~n1779 & ~n1788;
  assign n1794 = ~n1792 & n1793;
  assign n1795 = pi013 & ~pi014;
  assign n1796 = pi012 & ~n1795;
  assign n1797 = n1705 & ~n1796;
  assign n1798 = ~pi012 & ~n1664;
  assign n1799 = n408 & n1798;
  assign n1800 = ~n1717 & ~n1723;
  assign n1801 = ~n1750 & ~n1751;
  assign n1802 = n1800 & n1801;
  assign n1803 = ~n1672 & ~n1676;
  assign n1804 = ~n1745 & ~n1797;
  assign n1805 = n1803 & n1804;
  assign n1806 = n1692 & n1802;
  assign n1807 = ~n1707 & n1714;
  assign n1808 = n1721 & n1807;
  assign n1809 = n1805 & n1806;
  assign n1810 = ~n1695 & ~n1703;
  assign n1811 = n1762 & ~n1769;
  assign n1812 = ~n1774 & n1811;
  assign n1813 = n1809 & n1810;
  assign n1814 = ~n1666 & n1808;
  assign n1815 = ~n1756 & ~n1799;
  assign n1816 = n1814 & n1815;
  assign n1817 = n1812 & n1813;
  assign n1818 = n1794 & n1817;
  assign n1819 = n1816 & n1818;
  assign po014 = po020 | ~n1819;
  assign n1821 = ~po011 & ~po013;
  assign n1822 = ~po015 & n1821;
  assign po010 = po014 | ~n1822;
  assign n1824 = ~pi072 & ~pi074;
  assign n1825 = n1580 & ~n1824;
  assign n1826 = ~n368 & ~n442;
  assign n1827 = n622 & ~n1826;
  assign n1828 = n693 & n1669;
  assign n1829 = n438 & n1828;
  assign n1830 = ~pi010 & n1829;
  assign n1831 = n1660 & n1730;
  assign n1832 = ~n1665 & ~n1831;
  assign n1833 = ~n1830 & n1832;
  assign n1834 = n625 & n675;
  assign n1835 = n787 & n1834;
  assign n1836 = ~pi060 & n1835;
  assign n1837 = pi045 & n1836;
  assign n1838 = n1833 & ~n1837;
  assign n1839 = n492 & ~n1838;
  assign n1840 = ~n1029 & ~n1472;
  assign n1841 = n798 & ~n1840;
  assign n1842 = n664 & n1775;
  assign n1843 = n457 & n693;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = n465 & ~n1844;
  assign n1846 = ~n1841 & ~n1845;
  assign n1847 = n296 & ~n369;
  assign n1848 = ~n570 & ~n1847;
  assign n1849 = n416 & n740;
  assign n1850 = ~n1848 & n1849;
  assign n1851 = ~n434 & ~n1071;
  assign n1852 = n361 & ~n1851;
  assign n1853 = n1387 & n1852;
  assign n1854 = ~n1723 & ~n1853;
  assign n1855 = n630 & n1066;
  assign n1856 = n859 & n1718;
  assign n1857 = n507 & n599;
  assign n1858 = n376 & n510;
  assign n1859 = n1857 & n1858;
  assign n1860 = ~n1855 & ~n1856;
  assign n1861 = ~n1859 & n1860;
  assign n1862 = ~n1850 & n1854;
  assign n1863 = n1861 & n1862;
  assign n1864 = n1846 & n1863;
  assign n1865 = n419 & n1716;
  assign n1866 = ~n382 & ~n937;
  assign n1867 = n315 & ~n1866;
  assign n1868 = n315 & n616;
  assign n1869 = n1163 & n1868;
  assign n1870 = n315 & n508;
  assign n1871 = n1049 & n1870;
  assign n1872 = ~n1751 & ~n1871;
  assign n1873 = ~pi022 & n315;
  assign n1874 = ~pi021 & n420;
  assign n1875 = n1873 & n1874;
  assign n1876 = pi020 & n1875;
  assign n1877 = pi018 & n1876;
  assign n1878 = ~n1865 & ~n1869;
  assign n1879 = n1872 & n1878;
  assign n1880 = ~n1877 & n1879;
  assign n1881 = ~n1867 & n1880;
  assign n1882 = pi076 & ~n1881;
  assign n1883 = n312 & n369;
  assign n1884 = ~pi061 & n1513;
  assign n1885 = n798 & n1884;
  assign n1886 = n567 & n1102;
  assign n1887 = n573 & n1886;
  assign n1888 = ~n1885 & ~n1887;
  assign n1889 = n798 & n1345;
  assign n1890 = n1888 & ~n1889;
  assign n1891 = ~n1883 & n1890;
  assign n1892 = n308 & n744;
  assign n1893 = n349 & n1892;
  assign n1894 = ~n1138 & n1893;
  assign n1895 = n492 & n743;
  assign n1896 = n993 & n1895;
  assign n1897 = pi000 & n1896;
  assign n1898 = ~n1894 & ~n1897;
  assign n1899 = n1891 & n1898;
  assign n1900 = n480 & n971;
  assign n1901 = pi020 & n488;
  assign n1902 = ~n347 & ~n510;
  assign n1903 = n931 & ~n1902;
  assign n1904 = n354 & n508;
  assign n1905 = ~pi021 & n645;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = ~n1903 & n1906;
  assign n1908 = n293 & ~n1907;
  assign n1909 = ~n1900 & ~n1901;
  assign n1910 = ~n1908 & n1909;
  assign n1911 = ~n360 & ~n1910;
  assign n1912 = n471 & ~n1583;
  assign n1913 = pi060 & n1835;
  assign n1914 = n992 & n1892;
  assign n1915 = n1466 & n1914;
  assign n1916 = n717 & n1579;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n790 & n1917;
  assign n1919 = pi055 & pi056;
  assign n1920 = n454 & n761;
  assign n1921 = ~n1919 & n1920;
  assign n1922 = pi004 & pi006;
  assign n1923 = n781 & n1922;
  assign n1924 = ~n1913 & ~n1923;
  assign n1925 = ~n1921 & n1924;
  assign n1926 = ~n1226 & n1918;
  assign n1927 = n1925 & n1926;
  assign n1928 = n1912 & n1927;
  assign n1929 = n330 & ~n1928;
  assign n1930 = n454 & n1188;
  assign n1931 = n740 & n1930;
  assign n1932 = n667 & n1404;
  assign n1933 = n1243 & n1932;
  assign n1934 = n487 & n1076;
  assign n1935 = n354 & n509;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n1490 & n1936;
  assign n1938 = n938 & ~n1937;
  assign n1939 = pi011 & ~n1007;
  assign n1940 = pi013 & n1939;
  assign n1941 = ~n1718 & ~n1940;
  assign n1942 = n1368 & ~n1941;
  assign n1943 = n1485 & n1486;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1933 & n1944;
  assign n1946 = ~n1938 & n1945;
  assign n1947 = ~n1931 & n1946;
  assign n1948 = n335 & n549;
  assign n1949 = n311 & n1948;
  assign n1950 = n1217 & n1949;
  assign n1951 = n585 & n1950;
  assign n1952 = ~n1521 & ~n1915;
  assign n1953 = n1517 & ~n1952;
  assign n1954 = n369 & n416;
  assign n1955 = n334 & n1954;
  assign n1956 = ~n339 & ~n1955;
  assign n1957 = n1525 & ~n1956;
  assign n1958 = n1376 & n1521;
  assign n1959 = ~n1577 & ~n1951;
  assign n1960 = ~n1957 & n1959;
  assign n1961 = n1537 & n1960;
  assign n1962 = ~n1958 & n1961;
  assign n1963 = ~n1953 & n1962;
  assign n1964 = ~pi029 & n1304;
  assign n1965 = pi026 & n1964;
  assign n1966 = n1301 & n1965;
  assign n1967 = n477 & n479;
  assign n1968 = ~n360 & n1967;
  assign n1969 = n361 & n1366;
  assign n1970 = n417 & n1969;
  assign n1971 = pi007 & n1152;
  assign n1972 = ~pi001 & n1971;
  assign n1973 = ~n360 & n1972;
  assign n1974 = ~n1970 & ~n1973;
  assign n1975 = ~n360 & n593;
  assign n1976 = ~n363 & ~n1975;
  assign n1977 = n568 & ~n1976;
  assign n1978 = ~n1968 & n1974;
  assign n1979 = ~n1977 & n1978;
  assign n1980 = n740 & n1029;
  assign n1981 = n368 & n377;
  assign n1982 = n519 & n1981;
  assign n1983 = ~n1980 & ~n1982;
  assign n1984 = ~n711 & ~n1749;
  assign n1985 = ~pi013 & ~n1984;
  assign n1986 = n302 & n1670;
  assign n1987 = n299 & n1986;
  assign n1988 = ~pi011 & n1987;
  assign n1989 = pi013 & n303;
  assign n1990 = n438 & n1697;
  assign n1991 = ~n1671 & ~n1990;
  assign n1992 = n1989 & ~n1991;
  assign n1993 = pi045 & n1913;
  assign n1994 = n416 & n520;
  assign n1995 = ~n1158 & n1200;
  assign n1996 = pi015 & n465;
  assign n1997 = n1752 & n1996;
  assign n1998 = n787 & n1997;
  assign n1999 = ~n1138 & n1998;
  assign n2000 = n309 & n518;
  assign n2001 = n480 & n1396;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = n551 & ~n2002;
  assign n2004 = pi004 & n335;
  assign n2005 = ~n1398 & n2004;
  assign n2006 = ~n307 & n2005;
  assign n2007 = ~n722 & n734;
  assign n2008 = ~pi001 & n1396;
  assign n2009 = n687 & n2008;
  assign n2010 = n1396 & n1922;
  assign n2011 = n369 & n2010;
  assign n2012 = ~n2009 & ~n2011;
  assign n2013 = ~pi003 & ~n2012;
  assign n2014 = ~n400 & ~n973;
  assign n2015 = n418 & ~n2014;
  assign n2016 = n1379 & n2015;
  assign n2017 = ~n1466 & n1914;
  assign n2018 = ~pi122 & ~n1139;
  assign n2019 = n1140 & n2018;
  assign n2020 = ~n2017 & ~n2019;
  assign n2021 = n410 & n416;
  assign n2022 = n315 & n630;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = n420 & ~n2023;
  assign n2025 = n335 & n404;
  assign n2026 = ~n761 & ~n2025;
  assign n2027 = n336 & ~n2026;
  assign n2028 = n376 & n1491;
  assign n2029 = ~pi012 & n653;
  assign n2030 = ~pi013 & ~n580;
  assign n2031 = ~n2029 & n2030;
  assign n2032 = ~n1668 & ~n2031;
  assign n2033 = n460 & ~n2032;
  assign n2034 = n903 & ~n1450;
  assign n2035 = n1189 & n1401;
  assign n2036 = n798 & n2035;
  assign n2037 = pi122 & n1919;
  assign n2038 = n2036 & ~n2037;
  assign n2039 = n1228 & n1513;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = n427 & n1080;
  assign n2042 = n630 & n2041;
  assign n2043 = ~n1456 & ~n2042;
  assign n2044 = n904 & n1452;
  assign n2045 = n609 & n1670;
  assign n2046 = n585 & n2045;
  assign n2047 = n448 & n1990;
  assign n2048 = ~n290 & ~n607;
  assign n2049 = pi007 & ~n1783;
  assign n2050 = ~n2048 & n2049;
  assign n2051 = n442 & n2050;
  assign n2052 = n1787 & n2051;
  assign n2053 = n330 & n345;
  assign n2054 = n1435 & n2053;
  assign n2055 = pi011 & pi014;
  assign n2056 = ~pi013 & n1759;
  assign n2057 = ~n2055 & n2056;
  assign n2058 = n456 & n785;
  assign n2059 = ~pi009 & n625;
  assign n2060 = n2058 & n2059;
  assign n2061 = n302 & n607;
  assign n2062 = n2058 & n2061;
  assign n2063 = pi011 & n2062;
  assign n2064 = ~n2060 & ~n2063;
  assign n2065 = ~n2057 & n2064;
  assign n2066 = pi006 & ~n518;
  assign n2067 = ~pi007 & n2066;
  assign n2068 = n554 & n2067;
  assign n2069 = ~n2054 & ~n2068;
  assign n2070 = n2065 & n2069;
  assign n2071 = ~pi045 & n1836;
  assign n2072 = n798 & n2071;
  assign n2073 = ~n1138 & n1145;
  assign n2074 = ~pi021 & n436;
  assign n2075 = pi003 & n2008;
  assign n2076 = n549 & n2075;
  assign n2077 = pi020 & ~pi021;
  assign n2078 = n698 & n2077;
  assign n2079 = n320 & n589;
  assign n2080 = pi014 & n320;
  assign n2081 = n493 & n2080;
  assign n2082 = ~n2079 & ~n2081;
  assign n2083 = n635 & n2082;
  assign n2084 = ~n2078 & n2083;
  assign n2085 = n884 & n1161;
  assign n2086 = ~n360 & n528;
  assign n2087 = n596 & n1677;
  assign n2088 = n334 & n2087;
  assign n2089 = n428 & n2088;
  assign n2090 = ~n2086 & ~n2089;
  assign n2091 = pi001 & ~n2090;
  assign n2092 = n592 & n1715;
  assign n2093 = n1523 & n2092;
  assign n2094 = n330 & n1571;
  assign n2095 = ~n1133 & ~n2094;
  assign n2096 = n492 & n1463;
  assign n2097 = ~pi004 & ~pi006;
  assign n2098 = n555 & n2097;
  assign n2099 = n329 & ~n750;
  assign n2100 = n529 & n2010;
  assign n2101 = n404 & n1954;
  assign n2102 = ~n1225 & ~n1571;
  assign n2103 = n1234 & ~n2102;
  assign n2104 = ~n1139 & n1143;
  assign n2105 = ~pi122 & n2104;
  assign n2106 = ~n1207 & ~n2105;
  assign n2107 = ~n2103 & n2106;
  assign n2108 = ~pi022 & n1338;
  assign n2109 = n1313 & n2108;
  assign n2110 = n938 & n1243;
  assign n2111 = n699 & n2110;
  assign n2112 = n336 & n443;
  assign n2113 = ~n726 & ~n2112;
  assign n2114 = ~pi014 & n320;
  assign n2115 = n2113 & ~n2114;
  assign n2116 = ~n439 & n2115;
  assign n2117 = n332 & ~n2116;
  assign n2118 = ~n2100 & ~n2101;
  assign n2119 = ~n1994 & n2118;
  assign n2120 = ~n2003 & ~n2076;
  assign n2121 = ~n2098 & n2120;
  assign n2122 = ~n724 & n2119;
  assign n2123 = ~n1995 & ~n2006;
  assign n2124 = ~n2013 & ~n2016;
  assign n2125 = n2123 & n2124;
  assign n2126 = n2121 & n2122;
  assign n2127 = ~n1988 & ~n1999;
  assign n2128 = ~n2007 & ~n2024;
  assign n2129 = ~n2027 & ~n2085;
  assign n2130 = ~n2091 & ~n2099;
  assign n2131 = n2129 & n2130;
  assign n2132 = n2127 & n2128;
  assign n2133 = n2125 & n2126;
  assign n2134 = ~n1827 & ~n1993;
  assign n2135 = n2020 & n2040;
  assign n2136 = ~n2046 & ~n2047;
  assign n2137 = ~n2074 & ~n2093;
  assign n2138 = n2095 & ~n2096;
  assign n2139 = ~n2111 & n2138;
  assign n2140 = n2136 & n2137;
  assign n2141 = n2134 & n2135;
  assign n2142 = n2132 & n2133;
  assign n2143 = ~n1429 & n2131;
  assign n2144 = ~n1992 & ~n2028;
  assign n2145 = ~n2033 & ~n2034;
  assign n2146 = n2043 & ~n2052;
  assign n2147 = ~n2072 & ~n2073;
  assign n2148 = ~n2117 & n2147;
  assign n2149 = n2145 & n2146;
  assign n2150 = n2143 & n2144;
  assign n2151 = n2141 & n2142;
  assign n2152 = n2139 & n2140;
  assign n2153 = ~n1985 & ~n2044;
  assign n2154 = n2070 & n2084;
  assign n2155 = n2107 & ~n2109;
  assign n2156 = n2154 & n2155;
  assign n2157 = n2152 & n2153;
  assign n2158 = n2150 & n2151;
  assign n2159 = n2148 & n2149;
  assign n2160 = n696 & ~n1966;
  assign n2161 = n1979 & n1983;
  assign n2162 = n2160 & n2161;
  assign n2163 = n2158 & n2159;
  assign n2164 = n2156 & n2157;
  assign n2165 = n1794 & ~n1929;
  assign n2166 = n1947 & n1963;
  assign n2167 = n2165 & n2166;
  assign n2168 = n2163 & n2164;
  assign n2169 = n941 & n2162;
  assign n2170 = ~n1882 & n1899;
  assign n2171 = ~n1911 & n2170;
  assign n2172 = n2168 & n2169;
  assign n2173 = ~n1839 & n2167;
  assign n2174 = n1864 & n2173;
  assign n2175 = n2171 & n2172;
  assign n2176 = n2174 & n2175;
  assign n2177 = ~n1825 & n2176;
  assign n2178 = pi010 & n1731;
  assign n2179 = ~n1725 & ~n1997;
  assign n2180 = n1254 & ~n2179;
  assign n2181 = ~n2178 & ~n2180;
  assign n2182 = ~n368 & ~n1525;
  assign n2183 = n373 & ~n2182;
  assign n2184 = ~n1651 & ~n1737;
  assign n2185 = pi093 & n1649;
  assign n2186 = pi095 & n1735;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = n2184 & n2187;
  assign n2189 = ~n783 & n1093;
  assign n2190 = ~pi027 & n2189;
  assign n2191 = ~n1618 & ~n1628;
  assign n2192 = n492 & ~n2191;
  assign n2193 = ~n807 & n1627;
  assign n2194 = n492 & ~n2193;
  assign n2195 = n505 & ~n2194;
  assign n2196 = ~n2192 & n2195;
  assign po019 = n2190 | ~n2196;
  assign n2198 = pi005 & pi015;
  assign n2199 = n1641 & ~n2198;
  assign n2200 = ~pi012 & ~n1729;
  assign n2201 = n823 & ~n2200;
  assign n2202 = ~n589 & n2201;
  assign n2203 = ~n1644 & ~n2183;
  assign n2204 = ~n2199 & ~n2202;
  assign n2205 = n2203 & n2204;
  assign n2206 = ~n1727 & n2205;
  assign n2207 = ~n1653 & n2206;
  assign n2208 = ~n1739 & n2181;
  assign n2209 = n2207 & n2208;
  assign n2210 = ~po019 & n2209;
  assign n2211 = n2188 & n2210;
  assign po016 = ~n2177 | ~n2211;
  assign n2213 = n1011 & n1255;
  assign n2214 = n1306 & n1652;
  assign n2215 = pi009 & n2178;
  assign n2216 = ~n374 & ~n2201;
  assign n2217 = ~n2214 & n2216;
  assign n2218 = ~n2215 & n2217;
  assign n2219 = ~n2185 & ~n2213;
  assign n2220 = n2218 & n2219;
  assign po017 = ~n2177 | ~n2220;
  assign n2222 = ~n2186 & n2218;
  assign po018 = ~n2176 | ~n2222;
  assign n2224 = n346 & ~n1078;
  assign n2225 = n352 & n973;
  assign n2226 = n566 & n2225;
  assign n2227 = n1081 & n1365;
  assign n2228 = ~n2226 & ~n2227;
  assign n2229 = n776 & n1295;
  assign n2230 = ~n1275 & ~n1392;
  assign n2231 = n2228 & ~n2229;
  assign n2232 = n2230 & n2231;
  assign n2233 = n376 & n482;
  assign n2234 = ~n360 & n2233;
  assign n2235 = ~n2232 & n2234;
  assign n2236 = n1228 & n1472;
  assign n2237 = ~n1271 & ~n2236;
  assign n2238 = ~n1972 & n2237;
  assign n2239 = ~n360 & ~n2238;
  assign n2240 = ~n792 & ~n2239;
  assign n2241 = ~n487 & ~n1049;
  assign n2242 = n515 & ~n2241;
  assign n2243 = n354 & n484;
  assign n2244 = ~pi020 & n2243;
  assign n2245 = ~n2242 & ~n2244;
  assign n2246 = n1242 & n1243;
  assign n2247 = n1507 & ~n2246;
  assign n2248 = ~n794 & n2247;
  assign n2249 = n2245 & n2248;
  assign n2250 = ~n474 & ~n2249;
  assign n2251 = pi019 & n510;
  assign n2252 = ~n1527 & ~n2251;
  assign n2253 = n950 & ~n2252;
  assign n2254 = ~n384 & ~n410;
  assign n2255 = n1366 & ~n2254;
  assign n2256 = pi019 & n569;
  assign n2257 = ~n1259 & ~n2256;
  assign n2258 = n347 & n931;
  assign n2259 = n2257 & ~n2258;
  assign n2260 = ~n2255 & n2259;
  assign n2261 = n361 & ~n2260;
  assign n2262 = ~n1933 & ~n2261;
  assign n2263 = n1397 & n1922;
  assign n2264 = n480 & n550;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = n529 & ~n2265;
  assign n2267 = ~n937 & ~n1267;
  assign n2268 = ~n431 & ~n642;
  assign n2269 = n507 & ~n2268;
  assign n2270 = n354 & n2269;
  assign n2271 = n1492 & ~n2270;
  assign n2272 = n2267 & n2271;
  assign n2273 = n938 & ~n2272;
  assign n2274 = n514 & n1682;
  assign n2275 = n1069 & n1387;
  assign n2276 = ~pi022 & n2275;
  assign n2277 = ~n2274 & ~n2276;
  assign n2278 = n361 & ~n2277;
  assign n2279 = ~n1902 & n2229;
  assign n2280 = ~n592 & ~n1590;
  assign n2281 = n972 & ~n2280;
  assign n2282 = ~n2279 & ~n2281;
  assign n2283 = n938 & ~n2282;
  assign n2284 = ~n302 & ~n368;
  assign n2285 = n373 & ~n2284;
  assign n2286 = n518 & n1396;
  assign n2287 = ~n474 & n475;
  assign n2288 = n2286 & n2287;
  assign n2289 = n320 & n368;
  assign n2290 = n309 & n1170;
  assign n2291 = n480 & n2290;
  assign n2292 = ~n1393 & ~n2291;
  assign n2293 = ~n360 & ~n2292;
  assign n2294 = ~n416 & ~n453;
  assign n2295 = n552 & ~n2294;
  assign n2296 = pi001 & n454;
  assign n2297 = n310 & n2296;
  assign n2298 = ~n360 & n2297;
  assign n2299 = ~pi003 & n2298;
  assign n2300 = n518 & n719;
  assign n2301 = n376 & n1396;
  assign n2302 = n970 & n2301;
  assign n2303 = n345 & n2302;
  assign n2304 = ~n640 & ~n1103;
  assign n2305 = n345 & ~n2304;
  assign n2306 = ~n645 & ~n1102;
  assign n2307 = ~n356 & n2306;
  assign n2308 = n646 & ~n2307;
  assign n2309 = ~n2305 & ~n2308;
  assign po123 = n773 & n1161;
  assign n2311 = ~n1859 & ~po123;
  assign n2312 = ~n1279 & ~n1520;
  assign n2313 = ~pi039 & n360;
  assign n2314 = n1351 & ~n2313;
  assign n2315 = ~n1359 & ~n2314;
  assign n2316 = n2312 & n2315;
  assign n2317 = ~n1471 & n2316;
  assign n2318 = n330 & n797;
  assign n2319 = ~n596 & ~n630;
  assign n2320 = n2041 & ~n2319;
  assign n2321 = ~n2085 & ~n2320;
  assign n2322 = ~n2318 & n2321;
  assign n2323 = pi001 & n2301;
  assign n2324 = ~n392 & ~n2323;
  assign n2325 = ~pi122 & ~n2324;
  assign n2326 = n957 & n1397;
  assign n2327 = n992 & n2326;
  assign n2328 = ~n379 & ~n2327;
  assign n2329 = pi004 & n1397;
  assign n2330 = n349 & n2329;
  assign n2331 = n345 & n2330;
  assign n2332 = n1128 & n1397;
  assign n2333 = ~n381 & n2332;
  assign n2334 = n1396 & n1402;
  assign n2335 = n518 & n1397;
  assign n2336 = n992 & n2335;
  assign n2337 = ~n957 & ~n2097;
  assign n2338 = ~n360 & ~n2337;
  assign n2339 = n476 & n2338;
  assign n2340 = n528 & n551;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = ~n558 & ~n936;
  assign n2343 = ~n360 & n638;
  assign n2344 = n1516 & n2343;
  assign n2345 = ~n2333 & ~n2334;
  assign n2346 = ~n2336 & n2345;
  assign n2347 = ~n2325 & n2328;
  assign n2348 = ~n2331 & n2341;
  assign n2349 = n2347 & n2348;
  assign n2350 = n2346 & n2349;
  assign n2351 = ~n2344 & n2350;
  assign n2352 = n2322 & n2342;
  assign n2353 = n2351 & n2352;
  assign n2354 = ~n396 & n2353;
  assign n2355 = n972 & n1241;
  assign n2356 = n1243 & n2355;
  assign n2357 = ~pi057 & n2356;
  assign n2358 = n330 & n2357;
  assign n2359 = n359 & ~n1902;
  assign n2360 = n593 & n2359;
  assign n2361 = ~n2358 & ~n2360;
  assign n2362 = ~pi045 & ~n2361;
  assign n2363 = ~n1885 & n2040;
  assign n2364 = n1380 & n2021;
  assign n2365 = ~pi029 & ~pi045;
  assign n2366 = n568 & n2092;
  assign n2367 = ~pi082 & n2366;
  assign n2368 = n329 & n2367;
  assign n2369 = n2365 & n2368;
  assign n2370 = pi057 & n2356;
  assign n2371 = pi082 & n2366;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = n518 & n520;
  assign n2374 = n1275 & n2355;
  assign n2375 = n1378 & ~n1681;
  assign n2376 = n930 & n2375;
  assign n2377 = ~n2374 & ~n2376;
  assign n2378 = ~n2373 & n2377;
  assign n2379 = n2372 & n2378;
  assign n2380 = ~pi045 & ~n2379;
  assign n2381 = ~pi045 & n416;
  assign n2382 = n421 & n2381;
  assign n2383 = ~n2369 & ~n2382;
  assign n2384 = ~n2380 & n2383;
  assign n2385 = n2363 & ~n2364;
  assign n2386 = ~n2362 & n2385;
  assign n2387 = n2384 & n2386;
  assign n2388 = n1380 & n1868;
  assign n2389 = ~n1377 & n2388;
  assign n2390 = ~n580 & ~n653;
  assign n2391 = ~n302 & ~n2390;
  assign n2392 = ~n1728 & ~n2391;
  assign n2393 = n788 & ~n2392;
  assign n2394 = ~pi007 & n1485;
  assign n2395 = n336 & n2394;
  assign n2396 = n308 & n1485;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = ~n2393 & n2397;
  assign n2399 = ~n360 & ~n2398;
  assign n2400 = ~n2389 & ~n2399;
  assign n2401 = n1260 & n1763;
  assign n2402 = n1258 & n2401;
  assign n2403 = ~n1062 & ~n2402;
  assign n2404 = n506 & n717;
  assign n2405 = ~n348 & ~n2077;
  assign n2406 = pi018 & ~n2405;
  assign n2407 = n1712 & n2406;
  assign n2408 = ~n330 & ~n1517;
  assign n2409 = n1915 & ~n2408;
  assign n2410 = ~n1522 & ~n2409;
  assign n2411 = n347 & n667;
  assign n2412 = n1764 & n2411;
  assign n2413 = ~n966 & ~n2080;
  assign n2414 = n965 & ~n2413;
  assign n2415 = ~pi019 & n1385;
  assign n2416 = n348 & n2415;
  assign n2417 = n1081 & n2416;
  assign n2418 = ~n1090 & ~n2288;
  assign n2419 = ~n2289 & ~n2295;
  assign n2420 = ~n2300 & ~n2303;
  assign n2421 = n2419 & n2420;
  assign n2422 = ~n1968 & n2418;
  assign n2423 = ~n2266 & ~n2299;
  assign n2424 = n2422 & n2423;
  assign n2425 = ~n436 & n2421;
  assign n2426 = ~n1048 & ~n1084;
  assign n2427 = ~n1536 & ~n2285;
  assign n2428 = ~n2414 & ~n2417;
  assign n2429 = n2427 & n2428;
  assign n2430 = n2425 & n2426;
  assign n2431 = ~n617 & n2424;
  assign n2432 = ~n886 & ~n969;
  assign n2433 = ~n1067 & ~n2253;
  assign n2434 = ~n2404 & ~n2407;
  assign n2435 = ~n2412 & n2434;
  assign n2436 = n2432 & n2433;
  assign n2437 = n2430 & n2431;
  assign n2438 = ~n605 & n2429;
  assign n2439 = n1714 & n1854;
  assign n2440 = ~n2224 & n2311;
  assign n2441 = n2403 & n2440;
  assign n2442 = n2438 & n2439;
  assign n2443 = n2436 & n2437;
  assign n2444 = n2084 & n2435;
  assign n2445 = ~n2283 & ~n2293;
  assign n2446 = n2400 & n2410;
  assign n2447 = n2445 & n2446;
  assign n2448 = n2443 & n2444;
  assign n2449 = n2441 & n2442;
  assign n2450 = n366 & ~n2235;
  assign n2451 = ~n2278 & n2309;
  assign n2452 = n2450 & n2451;
  assign n2453 = n2448 & n2449;
  assign n2454 = ~n2273 & n2447;
  assign n2455 = n2453 & n2454;
  assign n2456 = n2262 & n2452;
  assign n2457 = n2317 & n2354;
  assign n2458 = n2456 & n2457;
  assign n2459 = ~n2250 & n2455;
  assign n2460 = n2387 & n2459;
  assign n2461 = n1460 & n2458;
  assign n2462 = n2240 & n2461;
  assign po022 = ~n2460 | ~n2462;
  assign n2464 = ~n1445 & n2387;
  assign n2465 = ~n374 & n2311;
  assign n2466 = n2322 & n2465;
  assign po023 = ~n2464 | ~n2466;
  assign n2468 = ~n360 & ~n2237;
  assign n2469 = ~n360 & ~n2247;
  assign n2470 = ~n1269 & ~n2469;
  assign n2471 = ~n360 & n1353;
  assign n2472 = ~n1440 & n1465;
  assign n2473 = n1376 & ~n2472;
  assign n2474 = ~pi021 & n1495;
  assign n2475 = n361 & n2394;
  assign n2476 = n1422 & ~n2475;
  assign n2477 = ~n2471 & ~n2474;
  assign n2478 = n2476 & n2477;
  assign n2479 = n2316 & ~n2473;
  assign n2480 = n2478 & n2479;
  assign n2481 = ~n2468 & n2480;
  assign n2482 = n2470 & n2481;
  assign po024 = ~n1413 | ~n2482;
  assign n2484 = n1424 & n1428;
  assign po025 = n1528 | n2484;
  assign n2486 = ~n1829 & n1832;
  assign n2487 = n437 & n1670;
  assign n2488 = ~n853 & ~n2487;
  assign n2489 = n585 & ~n2488;
  assign n2490 = n2486 & ~n2489;
  assign n2491 = n492 & ~n2490;
  assign n2492 = n692 & n1754;
  assign n2493 = ~n2491 & ~n2492;
  assign n2494 = n1080 & n1162;
  assign n2495 = n1244 & n2233;
  assign n2496 = ~pi020 & n2495;
  assign n2497 = ~n508 & ~n1371;
  assign n2498 = n1365 & ~n2497;
  assign n2499 = n1763 & n2498;
  assign n2500 = ~n2496 & ~n2499;
  assign n2501 = ~n1859 & n2500;
  assign n2502 = ~n2494 & n2501;
  assign n2503 = ~pi077 & ~n1692;
  assign n2504 = n519 & n1128;
  assign n2505 = n335 & n1397;
  assign n2506 = ~pi004 & n2505;
  assign n2507 = pi004 & ~pi006;
  assign n2508 = n525 & n2507;
  assign n2509 = ~n2506 & ~n2508;
  assign n2510 = pi005 & ~n2509;
  assign n2511 = n315 & n347;
  assign n2512 = pi018 & n2511;
  assign n2513 = n667 & n1276;
  assign n2514 = ~n2512 & ~n2513;
  assign n2515 = n487 & ~n2514;
  assign n2516 = n672 & n707;
  assign n2517 = pi012 & n1705;
  assign n2518 = n338 & n550;
  assign n2519 = n370 & n1396;
  assign po072 = n2518 | n2519;
  assign n2521 = n300 & n1669;
  assign n2522 = pi010 & n2521;
  assign n2523 = n898 & n2522;
  assign n2524 = ~n1987 & ~n2056;
  assign n2525 = ~pi011 & ~n2524;
  assign n2526 = ~n2523 & ~n2525;
  assign n2527 = ~po072 & n2526;
  assign n2528 = pi018 & n1766;
  assign n2529 = pi007 & pi010;
  assign n2530 = n300 & n2529;
  assign n2531 = ~pi009 & n2530;
  assign n2532 = n332 & n2531;
  assign n2533 = ~n2528 & ~n2532;
  assign n2534 = pi123 & ~n2533;
  assign n2535 = n852 & n2521;
  assign n2536 = ~pi010 & n2535;
  assign n2537 = ~n2534 & ~n2536;
  assign n2538 = pi020 & n1504;
  assign n2539 = pi020 & n1500;
  assign n2540 = n1228 & n2539;
  assign n2541 = pi018 & n2540;
  assign n2542 = ~n2538 & ~n2541;
  assign n2543 = n300 & n1780;
  assign n2544 = n494 & n2543;
  assign n2545 = n1418 & n2251;
  assign n2546 = n1385 & n2545;
  assign n2547 = ~n2332 & ~n2546;
  assign n2548 = pi007 & n299;
  assign n2549 = ~pi010 & n2548;
  assign n2550 = n609 & n1659;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = n898 & ~n2551;
  assign n2553 = n703 & n1671;
  assign n2554 = pi012 & n2553;
  assign n2555 = pi015 & n2554;
  assign n2556 = n1659 & n1718;
  assign n2557 = n299 & n2556;
  assign po115 = pi014 & n2557;
  assign n2559 = ~pi056 & ~pi080;
  assign n2560 = ~pi081 & ~pi082;
  assign n2561 = pi083 & n2560;
  assign n2562 = n2559 & n2561;
  assign n2563 = n1297 & n2562;
  assign n2564 = n510 & n2563;
  assign n2565 = ~pi065 & n2563;
  assign n2566 = n482 & n2565;
  assign n2567 = ~n2564 & ~n2566;
  assign n2568 = ~pi019 & n401;
  assign n2569 = pi022 & pi056;
  assign n2570 = n667 & n2569;
  assign n2571 = n376 & n2570;
  assign n2572 = n2568 & n2571;
  assign n2573 = n2567 & ~n2572;
  assign n2574 = n537 & ~n2573;
  assign n2575 = n1700 & n1728;
  assign n2576 = ~n1746 & n2575;
  assign n2577 = n789 & n1660;
  assign n2578 = n852 & n1990;
  assign n2579 = ~n1798 & ~n2578;
  assign n2580 = n854 & n1730;
  assign n2581 = ~n2577 & ~n2580;
  assign n2582 = n2579 & n2581;
  assign n2583 = n408 & ~n2582;
  assign n2584 = n408 & n1724;
  assign n2585 = ~n2488 & n2584;
  assign n2586 = ~n2576 & ~n2585;
  assign n2587 = ~n2583 & n2586;
  assign n2588 = ~n2574 & n2587;
  assign n2589 = pi061 & n2039;
  assign n2590 = n537 & n1294;
  assign n2591 = ~n2038 & ~n2590;
  assign n2592 = ~n2589 & n2591;
  assign n2593 = n2588 & n2592;
  assign n2594 = n580 & n1671;
  assign n2595 = pi012 & n2594;
  assign n2596 = n609 & n943;
  assign n2597 = n332 & n584;
  assign n2598 = n2596 & n2597;
  assign n2599 = ~n2046 & ~n2598;
  assign n2600 = ~pi014 & n332;
  assign n2601 = ~pi011 & n2600;
  assign n2602 = n2549 & n2601;
  assign n2603 = pi009 & n2602;
  assign n2604 = n2599 & ~n2603;
  assign n2605 = ~n2595 & n2604;
  assign n2606 = ~po115 & n2605;
  assign n2607 = n2593 & n2606;
  assign n2608 = ~n1216 & ~n1999;
  assign n2609 = n1236 & n2608;
  assign n2610 = n693 & n1789;
  assign n2611 = ~n409 & ~n1222;
  assign n2612 = ~n2610 & n2611;
  assign n2613 = n2609 & n2612;
  assign n2614 = ~n798 & ~n1338;
  assign n2615 = ~n330 & n2614;
  assign n2616 = ~n1315 & ~n2615;
  assign n2617 = ~n1966 & ~n2616;
  assign n2618 = pi035 & n492;
  assign n2619 = ~n799 & n1342;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = n1344 & ~n2620;
  assign n2622 = pi023 & n2621;
  assign n2623 = ~pi029 & n1753;
  assign n2624 = n2597 & n2623;
  assign n2625 = ~n2622 & ~n2624;
  assign n2626 = n2617 & n2625;
  assign n2627 = ~n2504 & ~n2510;
  assign n2628 = ~n2515 & ~n2516;
  assign n2629 = n2627 & n2628;
  assign n2630 = ~n2517 & ~n2544;
  assign n2631 = n2629 & n2630;
  assign n2632 = n2547 & ~n2552;
  assign n2633 = n2631 & n2632;
  assign n2634 = ~n2503 & ~n2555;
  assign n2635 = n2633 & n2634;
  assign n2636 = n2527 & n2542;
  assign n2637 = n2635 & n2636;
  assign n2638 = n2502 & n2537;
  assign n2639 = n2637 & n2638;
  assign n2640 = n2613 & n2639;
  assign n2641 = n2626 & n2640;
  assign n2642 = n2493 & n2641;
  assign po026 = ~n2607 | ~n2642;
  assign n2644 = ~pi026 & ~pi027;
  assign n2645 = ~pi045 & n2644;
  assign n2646 = n535 & n2645;
  assign n2647 = n1835 & n2646;
  assign n2648 = n1454 & ~n2647;
  assign n2649 = n1376 & n2539;
  assign n2650 = n2648 & ~n2649;
  assign n2651 = n653 & n1479;
  assign n2652 = n371 & n672;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = ~n1164 & n2653;
  assign n2655 = n596 & n1296;
  assign n2656 = n389 & n2655;
  assign n2657 = n2654 & ~n2656;
  assign n2658 = n345 & ~n2657;
  assign n2659 = ~n799 & n1436;
  assign n2660 = n511 & n1246;
  assign n2661 = n345 & n2660;
  assign n2662 = pi122 & ~n1919;
  assign n2663 = n492 & n2662;
  assign n2664 = ~n1455 & ~n2663;
  assign n2665 = n1435 & ~n2664;
  assign n2666 = ~n2659 & ~n2665;
  assign n2667 = ~n2661 & n2666;
  assign n2668 = pi020 & n2568;
  assign n2669 = n484 & n2668;
  assign n2670 = ~n1518 & n2669;
  assign n2671 = n1033 & n2080;
  assign n2672 = ~n1520 & ~n2671;
  assign n2673 = ~n2670 & n2672;
  assign n2674 = ~n360 & n740;
  assign n2675 = n1462 & n2674;
  assign n2676 = ~n1535 & ~n2675;
  assign n2677 = ~n344 & n492;
  assign n2678 = n1920 & n2677;
  assign n2679 = pi025 & n326;
  assign n2680 = n2644 & n2679;
  assign n2681 = ~n535 & ~n2680;
  assign n2682 = n1652 & ~n2681;
  assign n2683 = n1177 & ~n2294;
  assign n2684 = n518 & n1188;
  assign n2685 = pi007 & n2684;
  assign n2686 = ~n1294 & ~n2685;
  assign n2687 = ~n2683 & n2686;
  assign n2688 = n2677 & ~n2687;
  assign n2689 = ~n2053 & ~n2663;
  assign n2690 = n1177 & n1439;
  assign n2691 = ~n2689 & n2690;
  assign n2692 = pi028 & n739;
  assign n2693 = ~n328 & ~n2692;
  assign n2694 = ~n534 & ~n2693;
  assign n2695 = ~pi017 & n636;
  assign n2696 = n334 & n2695;
  assign n2697 = n377 & n2696;
  assign n2698 = n1036 & n2697;
  assign n2699 = ~n332 & n416;
  assign n2700 = n732 & n2699;
  assign n2701 = ~n2698 & ~n2700;
  assign n2702 = ~pi014 & n1955;
  assign n2703 = n1007 & n2702;
  assign n2704 = n291 & n963;
  assign n2705 = n300 & n2704;
  assign n2706 = n630 & n1582;
  assign n2707 = n1139 & n1142;
  assign n2708 = ~pi122 & n1620;
  assign n2709 = ~n503 & ~n2708;
  assign n2710 = n2707 & ~n2709;
  assign n2711 = ~n2705 & ~n2706;
  assign n2712 = ~n2710 & n2711;
  assign n2713 = n291 & n2597;
  assign n2714 = n299 & n2713;
  assign n2715 = n439 & n1674;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = pi012 & n2651;
  assign n2718 = ~pi122 & n2717;
  assign n2719 = n740 & n1501;
  assign n2720 = n359 & n1500;
  assign n2721 = n1517 & n2720;
  assign n2722 = ~n2719 & ~n2721;
  assign n2723 = ~n329 & ~n1228;
  assign n2724 = ~n360 & n1029;
  assign n2725 = ~n2723 & n2724;
  assign n2726 = n2722 & ~n2725;
  assign n2727 = ~n2694 & ~n2703;
  assign n2728 = ~n2678 & n2727;
  assign n2729 = ~n2691 & n2701;
  assign n2730 = n2728 & n2729;
  assign n2731 = n2676 & ~n2688;
  assign n2732 = n2730 & n2731;
  assign n2733 = ~n1279 & n2712;
  assign n2734 = n2716 & n2733;
  assign n2735 = n2673 & n2732;
  assign n2736 = ~n2682 & ~n2718;
  assign n2737 = n2735 & n2736;
  assign n2738 = n2667 & n2734;
  assign n2739 = n2737 & n2738;
  assign n2740 = ~n2658 & n2726;
  assign n2741 = n2739 & n2740;
  assign n2742 = n2650 & n2741;
  assign n2743 = ~pi122 & n329;
  assign n2744 = ~n2663 & ~n2743;
  assign n2745 = n1139 & n1143;
  assign n2746 = ~pi006 & n2745;
  assign n2747 = ~n2744 & n2746;
  assign n2748 = n1521 & n2053;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = ~n1953 & n2749;
  assign n2751 = n330 & ~n344;
  assign n2752 = n1309 & n2751;
  assign n2753 = pi029 & ~pi065;
  assign n2754 = n408 & ~n2753;
  assign n2755 = n1294 & n2754;
  assign n2756 = ~n1919 & n2755;
  assign n2757 = ~n2752 & ~n2756;
  assign n2758 = n1139 & n1140;
  assign n2759 = pi007 & n1440;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = n2663 & ~n2760;
  assign n2762 = n2757 & ~n2761;
  assign n2763 = ~pi029 & ~n360;
  assign n2764 = n416 & n2394;
  assign n2765 = n2763 & n2764;
  assign n2766 = n2762 & ~n2765;
  assign n2767 = n2750 & n2766;
  assign n2768 = n387 & n1049;
  assign n2769 = n484 & n2568;
  assign n2770 = ~n2768 & ~n2769;
  assign n2771 = ~pi018 & n1500;
  assign n2772 = n2770 & ~n2771;
  assign n2773 = ~n1328 & n2772;
  assign n2774 = n480 & n751;
  assign n2775 = n2773 & ~n2774;
  assign n2776 = n791 & ~n2775;
  assign n2777 = n416 & n1539;
  assign n2778 = n511 & n2777;
  assign n2779 = ~n2764 & ~n2778;
  assign n2780 = n438 & n1730;
  assign n2781 = n862 & n2780;
  assign n2782 = n2779 & ~n2781;
  assign n2783 = pi029 & ~n2782;
  assign n2784 = ~n2242 & n2324;
  assign n2785 = n507 & n1516;
  assign n2786 = ~n2244 & ~n2785;
  assign n2787 = n2784 & n2786;
  assign n2788 = ~pi122 & ~n2787;
  assign n2789 = pi088 & ~pi117;
  assign n2790 = n1527 & n2789;
  assign n2791 = n1352 & n2790;
  assign n2792 = n477 & n2789;
  assign n2793 = n315 & n2792;
  assign n2794 = ~n2791 & ~n2793;
  assign n2795 = ~n906 & n2794;
  assign n2796 = n329 & ~n2795;
  assign n2797 = pi023 & n592;
  assign n2798 = pi022 & n1870;
  assign n2799 = n2797 & n2798;
  assign n2800 = pi122 & n2799;
  assign n2801 = ~pi122 & n2246;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = n2311 & n2802;
  assign n2804 = ~n1326 & ~n2781;
  assign n2805 = ~pi029 & ~n2804;
  assign n2806 = ~n360 & n2805;
  assign n2807 = n2803 & ~n2806;
  assign n2808 = pi090 & n384;
  assign n2809 = n1579 & n2808;
  assign n2810 = pi092 & n384;
  assign n2811 = n1647 & n2810;
  assign n2812 = pi091 & n384;
  assign n2813 = n1646 & n2812;
  assign n2814 = ~pi096 & n1736;
  assign n2815 = n384 & ~n385;
  assign n2816 = n1648 & n2815;
  assign n2817 = ~n2814 & ~n2816;
  assign n2818 = ~pi097 & ~pi098;
  assign n2819 = ~n2817 & ~n2818;
  assign n2820 = ~n2811 & ~n2813;
  assign n2821 = n2188 & n2820;
  assign n2822 = ~n2819 & n2821;
  assign n2823 = ~n2809 & n2822;
  assign n2824 = ~n2285 & n2823;
  assign n2825 = n347 & n1857;
  assign n2826 = ~n297 & ~n2256;
  assign n2827 = ~n2825 & n2826;
  assign n2828 = ~n1886 & n2827;
  assign n2829 = n492 & ~n2828;
  assign n2830 = n938 & n2829;
  assign n2831 = ~pi029 & n511;
  assign n2832 = n327 & n737;
  assign n2833 = ~n738 & n2832;
  assign n2834 = ~n386 & ~n630;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = ~n2831 & ~n2835;
  assign n2837 = ~n360 & n2777;
  assign n2838 = ~n2836 & n2837;
  assign n2839 = n1325 & n1479;
  assign n2840 = n454 & n2394;
  assign n2841 = n465 & n1731;
  assign n2842 = ~n2839 & ~n2840;
  assign n2843 = ~n2841 & n2842;
  assign n2844 = ~n2833 & ~n2843;
  assign n2845 = ~pi020 & n347;
  assign n2846 = ~pi018 & n1243;
  assign n2847 = n2845 & n2846;
  assign n2848 = ~n2833 & n2847;
  assign n2849 = n416 & n2848;
  assign n2850 = ~n2844 & ~n2849;
  assign n2851 = ~n360 & ~n2850;
  assign n2852 = ~n2838 & ~n2851;
  assign n2853 = ~n1152 & ~n1892;
  assign n2854 = n349 & ~n2853;
  assign n2855 = ~n1215 & ~n1998;
  assign n2856 = ~n2854 & n2855;
  assign n2857 = ~n1186 & n2856;
  assign n2858 = n1151 & n2857;
  assign n2859 = ~n1138 & ~n2858;
  assign n2860 = ~n1146 & n1148;
  assign n2861 = n1202 & ~n1280;
  assign n2862 = ~n1194 & n2861;
  assign n2863 = ~n1221 & n2862;
  assign n2864 = ~n2860 & n2863;
  assign n2865 = ~n1158 & ~n2864;
  assign n2866 = ~n1196 & n2020;
  assign n2867 = n1184 & n2866;
  assign n2868 = n2107 & n2867;
  assign n2869 = ~n2865 & n2868;
  assign n2870 = ~n2859 & n2869;
  assign n2871 = ~n1896 & n2852;
  assign n2872 = n2870 & n2871;
  assign n2873 = n406 & n492;
  assign n2874 = ~n383 & ~n2873;
  assign n2875 = ~n393 & ~n2332;
  assign n2876 = ~n391 & n2875;
  assign n2877 = n2874 & n2876;
  assign n2878 = ~n381 & ~n2877;
  assign n2879 = n1163 & n2571;
  assign n2880 = pi065 & n2879;
  assign n2881 = n1376 & n2880;
  assign n2882 = n581 & n1255;
  assign n2883 = ~pi100 & n2882;
  assign n2884 = ~pi001 & ~n344;
  assign n2885 = pi122 & ~n2884;
  assign n2886 = n1971 & ~n2885;
  assign n2887 = n796 & ~n2886;
  assign n2888 = ~n2881 & n2887;
  assign n2889 = ~n2883 & n2888;
  assign n2890 = ~n2830 & n2889;
  assign n2891 = ~n2878 & n2890;
  assign n2892 = n2872 & n2891;
  assign n2893 = n1315 & ~n1345;
  assign n2894 = ~n2879 & n2893;
  assign n2895 = n791 & ~n2894;
  assign n2896 = ~n802 & ~n1095;
  assign n2897 = n1336 & ~n2896;
  assign n2898 = n789 & n1479;
  assign n2899 = ~n1883 & ~n2898;
  assign n2900 = ~n1920 & ~n2684;
  assign n2901 = n330 & ~n1919;
  assign n2902 = ~n2900 & n2901;
  assign n2903 = n492 & n961;
  assign n2904 = n963 & n2903;
  assign n2905 = n368 & ~n2413;
  assign n2906 = n929 & n930;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = ~n492 & ~n1376;
  assign n2909 = n1464 & ~n2908;
  assign n2910 = n606 & n944;
  assign n2911 = ~pi014 & n298;
  assign n2912 = n291 & n693;
  assign n2913 = n2911 & n2912;
  assign n2914 = ~pi008 & n2913;
  assign n2915 = n410 & n1638;
  assign n2916 = n1294 & n1965;
  assign n2917 = ~n344 & n2916;
  assign n2918 = n492 & n1916;
  assign n2919 = n771 & n1583;
  assign n2920 = ~pi122 & n2758;
  assign n2921 = ~n1915 & ~n2920;
  assign n2922 = n329 & ~n2921;
  assign n2923 = n1376 & n1463;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = n693 & n863;
  assign n2926 = ~n897 & ~n901;
  assign n2927 = n1724 & ~n2926;
  assign n2928 = ~n2925 & ~n2927;
  assign n2929 = ~n2093 & n2321;
  assign n2930 = n2928 & n2929;
  assign n2931 = ~n453 & ~n1922;
  assign n2932 = n970 & n1396;
  assign n2933 = ~n360 & n2932;
  assign n2934 = ~n2931 & n2933;
  assign n2935 = ~n1081 & ~n1418;
  assign n2936 = n1082 & ~n2935;
  assign n2937 = n361 & n2936;
  assign n2938 = n883 & n1539;
  assign n2939 = ~n599 & ~n1049;
  assign n2940 = n417 & ~n2939;
  assign n2941 = ~n2938 & ~n2940;
  assign n2942 = n1078 & n2941;
  assign n2943 = n346 & ~n2942;
  assign n2944 = pi012 & n725;
  assign n2945 = ~pi012 & n443;
  assign n2946 = ~n2944 & ~n2945;
  assign n2947 = ~pi015 & n308;
  assign n2948 = ~n2946 & n2947;
  assign n2949 = ~n1061 & ~n2948;
  assign n2950 = n359 & n2797;
  assign n2951 = ~n1857 & ~n2950;
  assign n2952 = ~n809 & n2951;
  assign n2953 = n928 & ~n2952;
  assign n2954 = ~n935 & n2949;
  assign n2955 = ~n2953 & n2954;
  assign n2956 = ~n2943 & n2955;
  assign n2957 = ~pi015 & n320;
  assign n2958 = n2600 & n2957;
  assign n2959 = ~n2253 & ~n2958;
  assign n2960 = ~n2339 & n2959;
  assign n2961 = n443 & n965;
  assign n2962 = ~n761 & ~n2961;
  assign n2963 = n314 & ~n2962;
  assign n2964 = n2083 & ~n2963;
  assign n2965 = ~n314 & ~n1922;
  assign n2966 = n719 & ~n2965;
  assign n2967 = n2960 & ~n2966;
  assign n2968 = n2964 & n2967;
  assign n2969 = ~n2937 & n2968;
  assign n2970 = n2956 & n2969;
  assign n2971 = n413 & n791;
  assign n2972 = ~n482 & n667;
  assign n2973 = ~n883 & ~n2972;
  assign n2974 = n1711 & ~n2973;
  assign n2975 = ~n362 & ~n773;
  assign n2976 = n1371 & ~n2975;
  assign n2977 = ~n1709 & ~n1722;
  assign n2978 = ~n2976 & n2977;
  assign n2979 = n376 & ~n2978;
  assign n2980 = ~n2974 & ~n2979;
  assign n2981 = ~n360 & ~n2980;
  assign n2982 = ~n2971 & ~n2981;
  assign n2983 = ~n2235 & n2982;
  assign n2984 = n2328 & n2983;
  assign n2985 = ~n2331 & ~n2934;
  assign n2986 = n2970 & n2985;
  assign n2987 = n2984 & n2986;
  assign n2988 = n1276 & n2846;
  assign n2989 = ~n2302 & ~n2988;
  assign n2990 = ~n2243 & n2989;
  assign n2991 = n345 & ~n2990;
  assign n2992 = ~n990 & n2035;
  assign n2993 = ~n344 & n2992;
  assign n2994 = n596 & n1246;
  assign n2995 = n2304 & ~n2994;
  assign n2996 = n1516 & n1680;
  assign n2997 = n2995 & ~n2996;
  assign n2998 = n345 & ~n2997;
  assign n2999 = pi023 & n2697;
  assign n3000 = n359 & n2999;
  assign n3001 = ~n2993 & ~n3000;
  assign n3002 = ~n2283 & n3001;
  assign n3003 = ~n2998 & n3002;
  assign n3004 = ~n2314 & ~n2991;
  assign n3005 = n3003 & n3004;
  assign n3006 = n2987 & n3005;
  assign n3007 = n329 & ~n820;
  assign n3008 = n329 & n405;
  assign n3009 = pi108 & pi109;
  assign n3010 = ~pi122 & n3009;
  assign n3011 = n827 & ~n3010;
  assign n3012 = n3008 & n3011;
  assign n3013 = ~n3007 & ~n3012;
  assign n3014 = pi029 & ~n3013;
  assign n3015 = ~n2318 & ~n3014;
  assign n3016 = pi022 & pi023;
  assign n3017 = n1284 & ~n3016;
  assign n3018 = n592 & n3017;
  assign n3019 = ~n1540 & ~n3018;
  assign n3020 = n1477 & n3019;
  assign n3021 = n416 & ~n3020;
  assign n3022 = n464 & n1255;
  assign n3023 = ~n1510 & ~n3022;
  assign n3024 = ~n1480 & ~n1482;
  assign n3025 = n3023 & n3024;
  assign n3026 = ~n1248 & ~n3021;
  assign n3027 = n3025 & n3026;
  assign n3028 = ~n1247 & n3027;
  assign n3029 = n1375 & ~n3028;
  assign n3030 = ~n2468 & ~n3029;
  assign n3031 = ~pi028 & ~n801;
  assign n3032 = ~n1262 & n1483;
  assign n3033 = n3031 & ~n3032;
  assign n3034 = n707 & n1718;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = ~n410 & ~n509;
  assign n3037 = n1065 & ~n3036;
  assign n3038 = n417 & n514;
  assign n3039 = n2306 & ~n3038;
  assign n3040 = ~n3037 & n3039;
  assign n3041 = n646 & ~n3040;
  assign n3042 = ~n2336 & ~n3041;
  assign n3043 = ~n360 & n1505;
  assign n3044 = n352 & n485;
  assign n3045 = n484 & n3044;
  assign n3046 = ~pi017 & n3045;
  assign n3047 = ~n2297 & ~n3046;
  assign n3048 = ~n1506 & n3047;
  assign n3049 = ~n360 & ~n3048;
  assign n3050 = ~n3043 & ~n3049;
  assign n3051 = ~n1727 & n2095;
  assign n3052 = n3050 & n3051;
  assign n3053 = n315 & n1523;
  assign n3054 = n1380 & n3053;
  assign n3055 = pi065 & n2564;
  assign n3056 = n1095 & n3055;
  assign n3057 = ~n1967 & ~n3056;
  assign n3058 = n520 & n1401;
  assign n3059 = n3057 & ~n3058;
  assign n3060 = ~n771 & ~n1228;
  assign n3061 = ~n2567 & ~n3060;
  assign n3062 = n771 & n2572;
  assign n3063 = ~n1431 & ~n3062;
  assign n3064 = ~n3061 & n3063;
  assign n3065 = n3059 & n3064;
  assign n3066 = ~n3054 & n3065;
  assign n3067 = ~n360 & ~n3066;
  assign n3068 = n385 & n930;
  assign n3069 = pi019 & n567;
  assign n3070 = ~n566 & n3069;
  assign n3071 = n1080 & n3070;
  assign n3072 = ~n3068 & ~n3071;
  assign n3073 = n293 & ~n3072;
  assign n3074 = n311 & ~n1358;
  assign n3075 = n1397 & ~n2931;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = n306 & ~n3076;
  assign n3078 = ~n3073 & ~n3077;
  assign n3079 = ~n360 & ~n3078;
  assign n3080 = n1071 & n3044;
  assign n3081 = n592 & n669;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = n598 & n1425;
  assign n3084 = ~n1902 & n3083;
  assign n3085 = ~n1902 & n2846;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = n3082 & n3086;
  assign n3088 = ~n511 & ~n596;
  assign n3089 = n353 & ~n3088;
  assign n3090 = n575 & n974;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = n3087 & n3091;
  assign n3093 = ~n1388 & ~n2255;
  assign n3094 = n2257 & n3093;
  assign n3095 = n3092 & n3094;
  assign n3096 = n361 & ~n3095;
  assign n3097 = n2400 & ~n3079;
  assign n3098 = ~n3096 & n3097;
  assign n3099 = n1148 & n1466;
  assign n3100 = ~n1462 & ~n3099;
  assign n3101 = ~n2689 & ~n3100;
  assign n3102 = n802 & n2662;
  assign n3103 = ~pi027 & ~n2693;
  assign n3104 = ~pi122 & n3103;
  assign n3105 = ~n2053 & ~n3102;
  assign n3106 = ~n3104 & n3105;
  assign n3107 = n1333 & ~n3106;
  assign n3108 = ~n3101 & ~n3107;
  assign n3109 = n693 & n897;
  assign n3110 = ~n1738 & ~n3109;
  assign n3111 = ~n330 & ~n791;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = ~n1440 & n3100;
  assign n3114 = n2743 & ~n3113;
  assign n3115 = n2053 & n2759;
  assign n3116 = n3108 & ~n3115;
  assign n3117 = ~n3112 & ~n3114;
  assign n3118 = n3116 & n3117;
  assign n3119 = ~n2914 & ~n2915;
  assign n3120 = ~n2917 & ~n2918;
  assign n3121 = ~n2919 & n3120;
  assign n3122 = ~n2902 & n3119;
  assign n3123 = ~n2910 & n3122;
  assign n3124 = n2899 & n3121;
  assign n3125 = ~n2904 & n2907;
  assign n3126 = ~n2909 & n3125;
  assign n3127 = n3123 & n3124;
  assign n3128 = n3126 & n3127;
  assign n3129 = n1233 & n1430;
  assign n3130 = ~n2788 & ~n2897;
  assign n3131 = n2924 & n2930;
  assign n3132 = n3130 & n3131;
  assign n3133 = n3128 & n3129;
  assign n3134 = ~n2273 & n2767;
  assign n3135 = ~n2776 & ~n2783;
  assign n3136 = n3042 & n3052;
  assign n3137 = n3135 & n3136;
  assign n3138 = n3133 & n3134;
  assign n3139 = ~n2796 & n3132;
  assign n3140 = n2807 & n3118;
  assign n3141 = n3139 & n3140;
  assign n3142 = n3137 & n3138;
  assign n3143 = ~n2895 & n3035;
  assign n3144 = n3098 & n3143;
  assign n3145 = n3141 & n3142;
  assign n3146 = n2464 & n2742;
  assign n3147 = ~n3067 & n3146;
  assign n3148 = n3144 & n3145;
  assign n3149 = n3015 & n3030;
  assign n3150 = n3148 & n3149;
  assign n3151 = n2892 & n3147;
  assign n3152 = n3006 & n3151;
  assign n3153 = n3150 & n3152;
  assign po027 = ~n2824 | ~n3153;
  assign n3155 = ~n1031 & ~n1572;
  assign n3156 = n1024 & ~n1939;
  assign n3157 = n713 & n1010;
  assign n3158 = n665 & ~n722;
  assign n3159 = ~n3156 & ~n3158;
  assign n3160 = n3155 & n3159;
  assign n3161 = n3157 & n3160;
  assign n3162 = n1101 & n3161;
  assign n3163 = n492 & n1219;
  assign n3164 = n798 & n1472;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = n676 & n963;
  assign n3167 = n2911 & n3166;
  assign n3168 = ~pi007 & n3167;
  assign n3169 = ~n717 & ~n1071;
  assign n3170 = n698 & ~n3169;
  assign n3171 = ~n1019 & ~n1053;
  assign n3172 = n751 & ~n3171;
  assign n3173 = ~n990 & n3172;
  assign n3174 = ~n1005 & ~n3173;
  assign n3175 = n1228 & n1571;
  assign n3176 = ~n344 & n3175;
  assign n3177 = ~pi015 & n728;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~n2224 & n3178;
  assign n3180 = n330 & n1336;
  assign n3181 = ~n1016 & ~n1026;
  assign n3182 = pi015 & ~n3181;
  assign n3183 = ~n990 & n1583;
  assign n3184 = ~n750 & ~n990;
  assign n3185 = ~n631 & ~n1044;
  assign n3186 = ~n3168 & ~n3183;
  assign n3187 = ~n3184 & n3186;
  assign n3188 = ~n1855 & n3185;
  assign n3189 = n3187 & n3188;
  assign n3190 = n1042 & ~n3170;
  assign n3191 = ~n3182 & n3190;
  assign n3192 = n3179 & n3189;
  assign n3193 = n3191 & n3192;
  assign n3194 = n2309 & ~n3180;
  assign n3195 = n3193 & n3194;
  assign n3196 = n3165 & n3195;
  assign n3197 = n3174 & n3196;
  assign n3198 = n565 & n3197;
  assign n3199 = n989 & n3198;
  assign po028 = ~n3162 | ~n3199;
  assign n3201 = ~n1785 & ~n2051;
  assign n3202 = n1673 & ~n3201;
  assign n3203 = pi031 & ~pi034;
  assign n3204 = ~n1597 & n3203;
  assign n3205 = ~n972 & n1625;
  assign n3206 = n429 & ~n3205;
  assign n3207 = ~pi127 & n455;
  assign n3208 = n338 & n375;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = ~pi002 & ~n3209;
  assign n3211 = n963 & n1950;
  assign n3212 = n425 & n2655;
  assign n3213 = n332 & n336;
  assign n3214 = n319 & n3213;
  assign n3215 = ~pi001 & n1397;
  assign n3216 = ~pi007 & n454;
  assign n3217 = n3215 & n3216;
  assign n3218 = ~n335 & ~n551;
  assign n3219 = n308 & n405;
  assign n3220 = ~n3218 & n3219;
  assign n3221 = ~pi004 & ~n453;
  assign n3222 = n730 & n3221;
  assign n3223 = n519 & n1948;
  assign n3224 = pi031 & pi034;
  assign n3225 = n1599 & ~n3224;
  assign n3226 = n751 & n1357;
  assign n3227 = pi007 & n611;
  assign n3228 = pi013 & ~n1007;
  assign n3229 = pi014 & n3228;
  assign n3230 = ~n584 & n3229;
  assign n3231 = n627 & n3230;
  assign n3232 = n628 & n1752;
  assign n3233 = pi021 & n1067;
  assign n3234 = n1834 & n2058;
  assign n3235 = ~n2062 & ~n3234;
  assign n3236 = ~pi029 & n869;
  assign n3237 = ~pi018 & n1504;
  assign n3238 = ~pi020 & n3237;
  assign n3239 = n680 & n2045;
  assign n3240 = n323 & n492;
  assign n3241 = pi014 & n676;
  assign n3242 = n1702 & n3241;
  assign n3243 = n1172 & n3242;
  assign n3244 = ~n732 & ~n3243;
  assign n3245 = n480 & ~n3244;
  assign n3246 = n823 & ~n1034;
  assign n3247 = n361 & n596;
  assign n3248 = pi020 & n1404;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = n487 & ~n3249;
  assign n3251 = n315 & n1387;
  assign n3252 = n386 & n3251;
  assign n3253 = ~n627 & ~n2522;
  assign n3254 = n450 & ~n3253;
  assign n3255 = ~n802 & ~n1376;
  assign n3256 = n1381 & ~n3255;
  assign n3257 = pi018 & ~pi029;
  assign n3258 = n329 & n3257;
  assign n3259 = n1500 & n3258;
  assign n3260 = n900 & n2780;
  assign n3261 = n416 & n482;
  assign n3262 = n2950 & n3261;
  assign n3263 = ~n3260 & ~n3262;
  assign n3264 = pi100 & n2882;
  assign n3265 = ~n581 & ~n1724;
  assign n3266 = n1754 & ~n3265;
  assign n3267 = ~pi023 & n510;
  assign n3268 = n315 & n566;
  assign n3269 = n773 & n3268;
  assign n3270 = n3267 & n3269;
  assign n3271 = ~n3266 & ~n3270;
  assign n3272 = ~n313 & ~n995;
  assign n3273 = ~n3172 & n3272;
  assign n3274 = ~pi020 & n2388;
  assign n3275 = n750 & ~n997;
  assign n3276 = pi001 & n311;
  assign n3277 = n480 & n3276;
  assign n3278 = ~pi007 & n3277;
  assign n3279 = n3273 & ~n3278;
  assign n3280 = n3275 & n3279;
  assign n3281 = ~n2357 & ~n3274;
  assign n3282 = n3280 & n3281;
  assign n3283 = n1002 & n3282;
  assign n3284 = n492 & ~n3283;
  assign n3285 = n368 & n622;
  assign n3286 = ~n571 & n1849;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n1285 & ~n1541;
  assign n3289 = ~n1253 & ~n3023;
  assign po048 = ~n3288 | n3289;
  assign n3291 = ~n1250 & ~po048;
  assign n3292 = n1264 & ~n3032;
  assign n3293 = n3291 & ~n3292;
  assign n3294 = n1228 & n2720;
  assign n3295 = n960 & n1697;
  assign n3296 = n1674 & n1746;
  assign n3297 = n3295 & n3296;
  assign n3298 = n1622 & ~n3297;
  assign n3299 = ~n3294 & n3298;
  assign n3300 = n898 & n2045;
  assign n3301 = n789 & n1670;
  assign n3302 = n300 & n3301;
  assign n3303 = ~n3300 & ~n3302;
  assign n3304 = ~n496 & n1918;
  assign n3305 = ~n2367 & n3304;
  assign n3306 = pi029 & ~n3305;
  assign n3307 = n1629 & n3303;
  assign n3308 = ~n3306 & n3307;
  assign n3309 = n329 & ~n3308;
  assign n3310 = ~n1754 & ~n3295;
  assign n3311 = n2597 & ~n3310;
  assign n3312 = ~pi013 & n580;
  assign n3313 = n1694 & n3312;
  assign n3314 = ~n3311 & ~n3313;
  assign n3315 = n465 & n785;
  assign n3316 = n702 & n3315;
  assign n3317 = n1949 & n3316;
  assign n3318 = ~n1126 & n1433;
  assign n3319 = ~pi006 & n1967;
  assign n3320 = ~n360 & n3319;
  assign n3321 = ~n1515 & ~n3317;
  assign n3322 = ~n3320 & n3321;
  assign n3323 = n3318 & n3322;
  assign n3324 = n1596 & ~n3203;
  assign n3325 = n492 & n763;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = ~pi124 & ~n3326;
  assign n3328 = n2614 & ~n2692;
  assign n3329 = n1029 & ~n3328;
  assign n3330 = pi015 & n448;
  assign n3331 = n492 & n3330;
  assign n3332 = ~n2488 & n3331;
  assign n3333 = n535 & ~n2645;
  assign n3334 = ~pi045 & n2680;
  assign n3335 = ~n3333 & ~n3334;
  assign po051 = n1836 & ~n3335;
  assign n3337 = pi021 & n778;
  assign n3338 = n1258 & n3337;
  assign n3339 = ~po051 & ~n3338;
  assign n3340 = ~n1982 & ~n3332;
  assign n3341 = n3339 & n3340;
  assign n3342 = ~n592 & ~n1366;
  assign n3343 = n972 & ~n3342;
  assign n3344 = ~n2279 & ~n3343;
  assign n3345 = n2271 & n3344;
  assign n3346 = n938 & ~n3345;
  assign n3347 = n438 & n2529;
  assign n3348 = n492 & n789;
  assign n3349 = n3347 & n3348;
  assign n3350 = n493 & n2050;
  assign n3351 = ~pi012 & n1784;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = n960 & ~n3352;
  assign n3354 = n2579 & ~n3353;
  assign n3355 = n492 & ~n3354;
  assign n3356 = n303 & n1790;
  assign n3357 = pi011 & ~n1746;
  assign n3358 = ~n494 & n3357;
  assign n3359 = n2623 & n3358;
  assign n3360 = ~n3349 & ~n3356;
  assign n3361 = ~n3359 & n3360;
  assign n3362 = ~n3355 & n3361;
  assign n3363 = n853 & n1776;
  assign n3364 = n330 & n3363;
  assign n3365 = n692 & n1700;
  assign n3366 = pi012 & pi014;
  assign n3367 = n584 & n2487;
  assign n3368 = n330 & n3367;
  assign n3369 = ~n3366 & n3368;
  assign n3370 = ~n3365 & ~n3369;
  assign n3371 = ~n3364 & n3370;
  assign n3372 = n1730 & n3347;
  assign n3373 = ~n1665 & ~n3372;
  assign n3374 = ~n1830 & n3373;
  assign n3375 = n330 & ~n3374;
  assign n3376 = n3371 & ~n3375;
  assign n3377 = n310 & ~n474;
  assign n3378 = n742 & n3377;
  assign n3379 = ~n493 & ~n589;
  assign n3380 = n320 & ~n3379;
  assign n3381 = n464 & n675;
  assign n3382 = n458 & n3381;
  assign n3383 = ~n3378 & ~n3380;
  assign n3384 = ~n3382 & n3383;
  assign n3385 = n2317 & n3384;
  assign n3386 = n1350 & n3385;
  assign n3387 = ~n3214 & ~n3223;
  assign n3388 = ~n3217 & n3387;
  assign n3389 = ~n3220 & ~n3222;
  assign n3390 = ~n3225 & n3389;
  assign n3391 = ~n3206 & n3388;
  assign n3392 = ~n3210 & ~n3211;
  assign n3393 = ~n3212 & ~n3226;
  assign n3394 = ~n3240 & ~n3246;
  assign n3395 = n3393 & n3394;
  assign n3396 = n3391 & n3392;
  assign n3397 = ~n1639 & n3390;
  assign n3398 = ~n3231 & n3235;
  assign n3399 = ~n3245 & ~n3250;
  assign n3400 = n3398 & n3399;
  assign n3401 = n3396 & n3397;
  assign n3402 = n1051 & n3395;
  assign n3403 = ~n1062 & n1645;
  assign n3404 = ~n1993 & ~n3202;
  assign n3405 = ~n3204 & ~n3227;
  assign n3406 = ~n3232 & ~n3239;
  assign n3407 = ~n3256 & ~n3259;
  assign n3408 = n3406 & n3407;
  assign n3409 = n3404 & n3405;
  assign n3410 = n3402 & n3403;
  assign n3411 = n3400 & n3401;
  assign n3412 = ~n1502 & n1634;
  assign n3413 = ~n2399 & ~n3233;
  assign n3414 = ~n3236 & ~n3252;
  assign n3415 = n3413 & n3414;
  assign n3416 = n3411 & n3412;
  assign n3417 = n3409 & n3410;
  assign n3418 = n2181 & n3408;
  assign n3419 = n2372 & ~n3238;
  assign n3420 = ~n3254 & n3263;
  assign n3421 = ~n3264 & n3287;
  assign n3422 = ~n3327 & ~n3329;
  assign n3423 = n3341 & n3422;
  assign n3424 = n3420 & n3421;
  assign n3425 = n3418 & n3419;
  assign n3426 = n3416 & n3417;
  assign n3427 = ~n2189 & n3415;
  assign n3428 = n3271 & n3427;
  assign n3429 = n3425 & n3426;
  assign n3430 = n3423 & n3424;
  assign n3431 = n1963 & ~n3284;
  assign n3432 = n3314 & ~n3346;
  assign n3433 = n3431 & n3432;
  assign n3434 = n3429 & n3430;
  assign n3435 = n1410 & n3428;
  assign n3436 = n2262 & n2470;
  assign n3437 = n3299 & ~n3309;
  assign n3438 = n3436 & n3437;
  assign n3439 = n3434 & n3435;
  assign n3440 = n1459 & n3433;
  assign n3441 = ~n2239 & n3293;
  assign n3442 = n3323 & n3362;
  assign n3443 = n3376 & n3442;
  assign n3444 = n3440 & n3441;
  assign n3445 = n3438 & n3439;
  assign n3446 = n3444 & n3445;
  assign n3447 = n1324 & n3443;
  assign n3448 = n3386 & n3447;
  assign po029 = ~n3446 | ~n3448;
  assign n3450 = ~pi123 & ~n2533;
  assign n3451 = n644 & n1242;
  assign n3452 = ~n1770 & ~n2530;
  assign n3453 = n852 & ~n3452;
  assign n3454 = n448 & n1770;
  assign n3455 = n308 & n2075;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = ~n2264 & ~n2326;
  assign n3458 = ~n2286 & n3457;
  assign n3459 = n335 & ~n3458;
  assign n3460 = n349 & n2001;
  assign n3461 = n345 & n3460;
  assign n3462 = n551 & n2286;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = n1712 & n2972;
  assign n3465 = pi004 & ~n530;
  assign n3466 = ~n453 & n3465;
  assign n3467 = ~pi003 & n307;
  assign n3468 = n369 & n3467;
  assign n3469 = ~n3466 & ~n3468;
  assign n3470 = n1396 & ~n3469;
  assign n3471 = n1366 & n1687;
  assign n3472 = n898 & n2550;
  assign n3473 = pi011 & n332;
  assign n3474 = n2550 & n3473;
  assign n3475 = ~n2557 & ~n3474;
  assign n3476 = pi014 & ~n1826;
  assign n3477 = ~n606 & ~n965;
  assign n3478 = ~n3476 & n3477;
  assign n3479 = n1749 & ~n3478;
  assign n3480 = n330 & n3353;
  assign n3481 = n384 & n2401;
  assign n3482 = pi020 & n3481;
  assign n3483 = ~n2327 & ~n2333;
  assign n3484 = n1170 & n2001;
  assign n3485 = ~pi122 & n3484;
  assign n3486 = n3483 & ~n3485;
  assign n3487 = n1011 & n2543;
  assign n3488 = n1787 & ~n3201;
  assign n3489 = n654 & n2521;
  assign n3490 = pi018 & n2495;
  assign n3491 = ~n1765 & ~n3490;
  assign n3492 = ~pi020 & ~n3491;
  assign n3493 = ~pi020 & n1709;
  assign n3494 = n359 & ~n567;
  assign n3495 = ~n1260 & n3494;
  assign n3496 = n362 & n3495;
  assign n3497 = ~n1261 & ~n3496;
  assign n3498 = ~n3493 & n3497;
  assign n3499 = n1385 & ~n3498;
  assign n3500 = ~n3451 & n3463;
  assign n3501 = ~n1686 & n3500;
  assign n3502 = ~n3459 & ~n3471;
  assign n3503 = ~n3479 & n3486;
  assign n3504 = n3502 & n3503;
  assign n3505 = ~n3464 & n3501;
  assign n3506 = ~n3470 & ~n3472;
  assign n3507 = ~n3480 & ~n3487;
  assign n3508 = ~n3489 & n3507;
  assign n3509 = n3505 & n3506;
  assign n3510 = ~n3453 & n3504;
  assign n3511 = n3456 & n3475;
  assign n3512 = ~n3482 & ~n3488;
  assign n3513 = n3511 & n3512;
  assign n3514 = n3509 & n3510;
  assign n3515 = n3508 & n3514;
  assign n3516 = ~n3450 & n3513;
  assign n3517 = ~n3492 & ~n3499;
  assign n3518 = n3516 & n3517;
  assign po030 = ~n3515 | ~n3518;
  assign n3520 = n308 & n2505;
  assign n3521 = n898 & n1759;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = n2527 & n3522;
  assign n3524 = n492 & n3363;
  assign n3525 = ~n2492 & ~n3524;
  assign n3526 = ~n2684 & ~n2880;
  assign n3527 = n740 & ~n3526;
  assign n3528 = ~n1501 & ~n1513;
  assign n3529 = n1228 & ~n3528;
  assign n3530 = n680 & ~n1746;
  assign n3531 = n1754 & n3530;
  assign n3532 = n451 & ~n2488;
  assign n3533 = pi029 & n3532;
  assign n3534 = ~n1695 & ~n3533;
  assign n3535 = ~n3531 & n3534;
  assign n3536 = n581 & n2623;
  assign n3537 = ~n2042 & n2311;
  assign n3538 = n2753 & n2879;
  assign n3539 = n329 & n3538;
  assign n3540 = n2486 & ~n3367;
  assign n3541 = n492 & ~n3540;
  assign n3542 = n330 & n3277;
  assign n3543 = n1076 & n2041;
  assign n3544 = ~pi020 & n330;
  assign n3545 = n1500 & n3544;
  assign n3546 = n2591 & ~n3545;
  assign n3547 = n2617 & n3546;
  assign n3548 = ~pi015 & n2603;
  assign n3549 = ~n1705 & ~n3542;
  assign n3550 = ~n3543 & n3549;
  assign n3551 = ~n2046 & ~n2553;
  assign n3552 = ~n2621 & n3551;
  assign n3553 = ~n2538 & n3550;
  assign n3554 = ~n3539 & n3553;
  assign n3555 = n1888 & n3552;
  assign n3556 = ~n3527 & ~n3529;
  assign n3557 = ~n3536 & n3537;
  assign n3558 = ~n3548 & n3557;
  assign n3559 = n3555 & n3556;
  assign n3560 = ~n1792 & n3554;
  assign n3561 = n3525 & n3560;
  assign n3562 = n3558 & n3559;
  assign n3563 = n2537 & n3523;
  assign n3564 = n3535 & n3563;
  assign n3565 = n3561 & n3562;
  assign n3566 = n3564 & n3565;
  assign n3567 = ~n3541 & n3547;
  assign n3568 = n3566 & n3567;
  assign po031 = ~n2588 | ~n3568;
  assign n3570 = pi017 & n1687;
  assign n3571 = n2225 & n3570;
  assign n3572 = ~n2358 & n2377;
  assign n3573 = n304 & n2522;
  assign n3574 = ~n3571 & ~n3573;
  assign n3575 = n3572 & n3574;
  assign n3576 = ~pi023 & ~n347;
  assign n3577 = ~n1365 & ~n3576;
  assign n3578 = n1684 & n3577;
  assign n3579 = n1295 & n3578;
  assign n3580 = ~pi023 & n315;
  assign n3581 = pi022 & ~n1708;
  assign n3582 = ~n883 & ~n3581;
  assign n3583 = n3580 & ~n3582;
  assign n3584 = pi018 & ~n347;
  assign n3585 = n1715 & n3584;
  assign n3586 = ~n3583 & ~n3585;
  assign n3587 = n644 & ~n3586;
  assign n3588 = ~n3579 & ~n3587;
  assign n3589 = n1872 & n3588;
  assign n3590 = n1378 & n1405;
  assign n3591 = n486 & n1684;
  assign n3592 = n1284 & n3591;
  assign n3593 = ~n3590 & ~n3592;
  assign n3594 = n717 & n1711;
  assign n3595 = ~pi013 & ~n3366;
  assign n3596 = n1749 & n3595;
  assign n3597 = n453 & n550;
  assign n3598 = n3465 & n3597;
  assign n3599 = n315 & n3083;
  assign n3600 = pi023 & n2511;
  assign n3601 = n1425 & n3600;
  assign n3602 = n774 & n3580;
  assign n3603 = n420 & n1870;
  assign n3604 = n507 & n1378;
  assign n3605 = n315 & n642;
  assign n3606 = n2077 & n3605;
  assign n3607 = ~pi018 & n3600;
  assign n3608 = ~n3604 & ~n3606;
  assign n3609 = ~n3607 & n3608;
  assign n3610 = n773 & ~n3609;
  assign n3611 = ~n3603 & ~n3610;
  assign n3612 = ~n3602 & n3611;
  assign n3613 = n315 & n1027;
  assign n3614 = n420 & n3613;
  assign n3615 = ~pi023 & n3614;
  assign n3616 = n3612 & ~n3615;
  assign n3617 = n420 & n667;
  assign n3618 = ~pi020 & n1539;
  assign n3619 = ~n2668 & ~n3618;
  assign n3620 = ~n3617 & n3619;
  assign n3621 = n354 & n566;
  assign n3622 = n3620 & ~n3621;
  assign n3623 = n2511 & ~n3622;
  assign n3624 = n1070 & n3591;
  assign n3625 = n3616 & ~n3624;
  assign n3626 = ~n3623 & n3625;
  assign n3627 = ~n3601 & n3626;
  assign n3628 = ~pi023 & n417;
  assign n3629 = n1685 & n3628;
  assign n3630 = ~n1723 & ~n3269;
  assign n3631 = ~n3629 & n3630;
  assign n3632 = ~pi022 & ~n3631;
  assign n3633 = ~n1377 & n3274;
  assign n3634 = n315 & n1527;
  assign n3635 = n1081 & n3634;
  assign n3636 = n1874 & n3268;
  assign n3637 = n630 & n1516;
  assign n3638 = n492 & n3637;
  assign n3639 = ~pi019 & ~pi021;
  assign n3640 = n1425 & n3639;
  assign n3641 = n1873 & n3640;
  assign n3642 = n1378 & n1681;
  assign n3643 = ~n3613 & ~n3642;
  assign n3644 = n487 & ~n3643;
  assign n3645 = n772 & n1716;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = ~n3636 & n3646;
  assign n3648 = ~n3641 & n3647;
  assign n3649 = ~n3638 & n3648;
  assign n3650 = n644 & n1688;
  assign n3651 = ~pi029 & n2368;
  assign n3652 = ~n1757 & ~n2009;
  assign n3653 = ~n3598 & ~n3650;
  assign n3654 = n3652 & n3653;
  assign n3655 = ~n2417 & ~n3594;
  assign n3656 = ~n3596 & ~n3635;
  assign n3657 = n3655 & n3656;
  assign n3658 = ~n2344 & n3654;
  assign n3659 = ~n3599 & n3658;
  assign n3660 = ~n1876 & n3657;
  assign n3661 = n3589 & ~n3633;
  assign n3662 = n3660 & n3661;
  assign n3663 = n3593 & n3659;
  assign n3664 = ~n3632 & n3663;
  assign n3665 = ~n1867 & n3662;
  assign n3666 = n3575 & n3649;
  assign n3667 = ~n3651 & n3666;
  assign n3668 = n3664 & n3665;
  assign n3669 = n3667 & n3668;
  assign po032 = ~n3627 | ~n3669;
  assign n3671 = n2301 & ~n3218;
  assign n3672 = n974 & n1242;
  assign n3673 = n789 & n2543;
  assign n3674 = ~n368 & ~n1752;
  assign n3675 = n1772 & ~n3674;
  assign n3676 = n1712 & n2845;
  assign n3677 = n290 & n606;
  assign n3678 = n609 & n3677;
  assign n3679 = ~pi007 & n3678;
  assign n3680 = n1366 & n1688;
  assign n3681 = n412 & n1385;
  assign n3682 = ~n1770 & ~n2596;
  assign n3683 = n2597 & ~n3682;
  assign n3684 = ~n3671 & ~n3672;
  assign n3685 = ~n3680 & n3684;
  assign n3686 = ~n3673 & ~n3675;
  assign n3687 = ~n3676 & ~n3679;
  assign n3688 = ~n3681 & n3687;
  assign n3689 = n3685 & n3686;
  assign n3690 = ~n3683 & n3689;
  assign po033 = ~n3688 | ~n3690;
  assign n3692 = n492 & n741;
  assign n3693 = pi124 & ~n3326;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = ~pi017 & n3212;
  assign n3696 = pi064 & n3695;
  assign n3697 = n429 & ~n1625;
  assign n3698 = n1595 & ~n3203;
  assign n3699 = ~n824 & ~n3223;
  assign n3700 = ~n3697 & n3699;
  assign n3701 = ~n3338 & ~n3698;
  assign n3702 = n3700 & n3701;
  assign n3703 = ~n3696 & n3702;
  assign po034 = ~n3694 | ~n3703;
  assign n3705 = n675 & n1842;
  assign n3706 = pi023 & n3233;
  assign n3707 = ~n2724 & n2921;
  assign n3708 = ~n1335 & n3707;
  assign n3709 = n818 & n828;
  assign n3710 = pi012 & n1661;
  assign n3711 = ~n1830 & ~n2367;
  assign n3712 = ~n3710 & n3711;
  assign n3713 = ~n3709 & n3712;
  assign n3714 = pi029 & ~n3713;
  assign n3715 = ~n468 & ~n797;
  assign n3716 = ~n814 & n3715;
  assign n3717 = n3708 & n3716;
  assign n3718 = ~n3714 & n3717;
  assign n3719 = n329 & ~n3718;
  assign n3720 = n938 & ~n2832;
  assign n3721 = n2847 & n3720;
  assign n3722 = ~n497 & ~n3721;
  assign n3723 = ~n574 & ~n1088;
  assign n3724 = ~n2783 & n3722;
  assign n3725 = n3723 & n3724;
  assign n3726 = n345 & n2652;
  assign n3727 = ~pi014 & n3726;
  assign n3728 = n492 & n2791;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = ~n2670 & n3729;
  assign n3731 = n589 & ~n2413;
  assign n3732 = n361 & n3085;
  assign n3733 = ~n2677 & ~n2901;
  assign n3734 = n1920 & ~n3733;
  assign n3735 = pi015 & n3734;
  assign n3736 = ~pi019 & n413;
  assign n3737 = ~n3109 & ~n3736;
  assign n3738 = n791 & ~n3737;
  assign n3739 = ~pi019 & n391;
  assign n3740 = ~n381 & n3739;
  assign n3741 = n1071 & n1975;
  assign n3742 = ~n3740 & ~n3741;
  assign n3743 = ~n477 & ~n2256;
  assign n3744 = n604 & ~n3743;
  assign n3745 = n928 & n2950;
  assign n3746 = n1426 & n1428;
  assign n3747 = pi019 & n3746;
  assign n3748 = ~n3735 & ~n3744;
  assign n3749 = ~n3745 & ~n3747;
  assign n3750 = n3748 & n3749;
  assign n3751 = n3742 & n3750;
  assign n3752 = ~n3738 & n3751;
  assign n3753 = ~n3731 & ~n3732;
  assign n3754 = n3730 & n3753;
  assign n3755 = n3752 & n3754;
  assign n3756 = n642 & n3337;
  assign n3757 = ~n360 & n483;
  assign n3758 = pi020 & n3757;
  assign n3759 = n1275 & n3758;
  assign n3760 = ~n3756 & ~n3759;
  assign n3761 = ~pi018 & ~n3760;
  assign n3762 = ~n1095 & ~n1569;
  assign n3763 = n1571 & ~n3762;
  assign n3764 = ~n591 & ~n3763;
  assign n3765 = ~n2958 & n3764;
  assign n3766 = n940 & n3765;
  assign n3767 = ~n3761 & n3766;
  assign n3768 = n802 & n1333;
  assign n3769 = ~n2037 & n3768;
  assign n3770 = ~pi011 & n1659;
  assign n3771 = pi012 & n3770;
  assign n3772 = n692 & n1697;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = n1673 & ~n3773;
  assign n3775 = n771 & ~n780;
  assign n3776 = n487 & n938;
  assign n3777 = ~n1066 & ~n3776;
  assign n3778 = n717 & ~n3777;
  assign n3779 = pi005 & n1640;
  assign n3780 = ~n824 & ~n3779;
  assign n3781 = pi015 & ~n3780;
  assign n3782 = ~n2690 & n2760;
  assign n3783 = n2663 & ~n3782;
  assign n3784 = pi108 & ~n1002;
  assign n3785 = n991 & ~n3784;
  assign n3786 = ~n828 & ~n990;
  assign n3787 = ~n3785 & n3786;
  assign n3788 = ~n328 & ~n537;
  assign n3789 = n532 & ~n3788;
  assign n3790 = ~n329 & n2614;
  assign n3791 = n533 & ~n3790;
  assign n3792 = ~n3789 & ~n3791;
  assign n3793 = ~pi089 & ~n587;
  assign n3794 = n582 & n620;
  assign n3795 = ~n586 & ~n3794;
  assign n3796 = ~n3793 & n3795;
  assign n3797 = ~pi012 & n345;
  assign n3798 = n2651 & n3797;
  assign n3799 = n3796 & ~n3798;
  assign n3800 = n3792 & n3799;
  assign n3801 = ~n3081 & ~n3090;
  assign n3802 = n410 & n598;
  assign n3803 = n389 & n3802;
  assign n3804 = n3801 & ~n3803;
  assign n3805 = ~n2258 & n3804;
  assign n3806 = n293 & ~n3805;
  assign n3807 = n788 & n1718;
  assign n3808 = n482 & n810;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = ~n3806 & n3809;
  assign n3811 = ~n474 & ~n3810;
  assign n3812 = n1262 & n3031;
  assign n3813 = n1064 & n2999;
  assign n3814 = n896 & n899;
  assign n3815 = ~n1583 & ~n3814;
  assign n3816 = n3103 & ~n3815;
  assign n3817 = ~n990 & ~n3275;
  assign n3818 = n329 & n470;
  assign n3819 = pi029 & pi067;
  assign n3820 = n3818 & ~n3819;
  assign n3821 = ~n2906 & ~n3813;
  assign n3822 = ~n3817 & n3821;
  assign n3823 = ~n3820 & n3822;
  assign n3824 = ~n3816 & n3823;
  assign n3825 = n832 & n3008;
  assign n3826 = n329 & n818;
  assign n3827 = ~n879 & ~n3826;
  assign n3828 = ~n816 & ~n3827;
  assign n3829 = n877 & ~n3825;
  assign n3830 = ~n3828 & n3829;
  assign n3831 = ~pi029 & n2682;
  assign n3832 = n896 & n904;
  assign n3833 = n740 & n3832;
  assign n3834 = n1336 & n2692;
  assign n3835 = ~n3831 & ~n3833;
  assign n3836 = ~n3834 & n3835;
  assign n3837 = n3165 & n3836;
  assign n3838 = n386 & n2777;
  assign n3839 = ~n2839 & ~n3838;
  assign n3840 = ~n474 & ~n2832;
  assign n3841 = ~n3839 & n3840;
  assign n3842 = n735 & n1033;
  assign n3843 = ~n828 & n3842;
  assign n3844 = ~n584 & ~n3530;
  assign n3845 = n460 & ~n3844;
  assign n3846 = ~n688 & ~n1089;
  assign n3847 = n319 & ~n3846;
  assign n3848 = ~n1032 & ~n3847;
  assign n3849 = ~pi015 & ~n3848;
  assign n3850 = ~pi010 & n692;
  assign n3851 = n664 & n3850;
  assign n3852 = n1006 & n1728;
  assign n3853 = n622 & n3852;
  assign n3854 = n938 & n1523;
  assign n3855 = n1366 & n3854;
  assign n3856 = n581 & n1753;
  assign n3857 = pi029 & n3856;
  assign n3858 = n332 & n734;
  assign n3859 = n621 & n692;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = pi014 & ~n3860;
  assign n3862 = n609 & n2713;
  assign n3863 = ~n2715 & ~n3862;
  assign n3864 = n646 & ~n2306;
  assign n3865 = n2097 & n2600;
  assign n3866 = n319 & n3865;
  assign n3867 = ~pi015 & n3866;
  assign n3868 = n345 & ~n2995;
  assign n3869 = ~pi113 & n1462;
  assign n3870 = ~n3099 & ~n3869;
  assign n3871 = ~n2037 & ~n3870;
  assign n3872 = ~pi122 & n1440;
  assign n3873 = ~n1916 & ~n3872;
  assign n3874 = ~n2388 & n3873;
  assign n3875 = ~n807 & ~n1464;
  assign n3876 = n3874 & n3875;
  assign n3877 = ~n3871 & n3876;
  assign n3878 = n492 & ~n3877;
  assign n3879 = ~n566 & ~n668;
  assign n3880 = n1428 & ~n3879;
  assign n3881 = n1590 & n3880;
  assign n3882 = ~n340 & ~n723;
  assign n3883 = n368 & ~n3882;
  assign n3884 = ~n508 & ~n511;
  assign n3885 = pi019 & ~n3884;
  assign n3886 = n363 & n3885;
  assign n3887 = n678 & n898;
  assign n3888 = ~n630 & ~n883;
  assign n3889 = pi023 & n429;
  assign n3890 = ~n3888 & n3889;
  assign n3891 = n827 & ~n834;
  assign n3892 = ~n831 & n3891;
  assign n3893 = n314 & n2961;
  assign n3894 = ~pi014 & n734;
  assign n3895 = n330 & n405;
  assign n3896 = n829 & n3895;
  assign n3897 = ~pi010 & n442;
  assign n3898 = n620 & n3897;
  assign n3899 = n2055 & n3898;
  assign n3900 = n1024 & ~n1728;
  assign n3901 = n791 & n2769;
  assign n3902 = pi023 & n578;
  assign n3903 = n599 & n2021;
  assign n3904 = ~n2360 & ~n3903;
  assign n3905 = n387 & n2568;
  assign n3906 = n408 & n3905;
  assign n3907 = n707 & n852;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = ~n711 & n3908;
  assign n3910 = ~pi011 & n1009;
  assign n3911 = ~n3902 & ~n3910;
  assign n3912 = ~n414 & n3911;
  assign n3913 = n3904 & n3912;
  assign n3914 = n3909 & n3913;
  assign n3915 = ~n3867 & ~n3881;
  assign n3916 = ~n3893 & ~n3896;
  assign n3917 = n3915 & n3916;
  assign n3918 = ~n662 & ~n2915;
  assign n3919 = ~n3843 & ~n3851;
  assign n3920 = ~n3855 & ~n3883;
  assign n3921 = ~n3886 & ~n3887;
  assign n3922 = ~n3890 & ~n3894;
  assign n3923 = ~n3899 & n3922;
  assign n3924 = n3920 & n3921;
  assign n3925 = n3918 & n3919;
  assign n3926 = ~n706 & n3917;
  assign n3927 = ~n3705 & ~n3774;
  assign n3928 = ~n3781 & ~n3849;
  assign n3929 = ~n3853 & ~n3892;
  assign n3930 = ~n3901 & n3929;
  assign n3931 = n3927 & n3928;
  assign n3932 = n3925 & n3926;
  assign n3933 = n3923 & n3924;
  assign n3934 = n1063 & ~n2371;
  assign n3935 = n2712 & ~n3294;
  assign n3936 = ~n3778 & ~n3845;
  assign n3937 = ~n3861 & n3863;
  assign n3938 = ~n3864 & ~n3900;
  assign n3939 = n3937 & n3938;
  assign n3940 = n3935 & n3936;
  assign n3941 = n3933 & n3934;
  assign n3942 = n3931 & n3932;
  assign n3943 = n1023 & n3930;
  assign n3944 = ~n1031 & n3179;
  assign n3945 = n3370 & ~n3706;
  assign n3946 = ~n3769 & ~n3775;
  assign n3947 = ~n3783 & ~n3812;
  assign n3948 = ~n3857 & n3947;
  assign n3949 = n3945 & n3946;
  assign n3950 = n3943 & n3944;
  assign n3951 = n3941 & n3942;
  assign n3952 = n3939 & n3940;
  assign n3953 = n463 & n1979;
  assign n3954 = n2750 & n3767;
  assign n3955 = ~n3841 & ~n3868;
  assign n3956 = n3954 & n3955;
  assign n3957 = n3952 & n3953;
  assign n3958 = n3950 & n3951;
  assign n3959 = n3948 & n3949;
  assign n3960 = n3314 & ~n3787;
  assign n3961 = n3824 & ~n3878;
  assign n3962 = n3914 & n3961;
  assign n3963 = n3959 & n3960;
  assign n3964 = n3957 & n3958;
  assign n3965 = n3800 & n3956;
  assign n3966 = ~n3811 & n3965;
  assign n3967 = n3963 & n3964;
  assign n3968 = n861 & n3962;
  assign n3969 = n3725 & n3755;
  assign n3970 = n3830 & n3837;
  assign n3971 = n3969 & n3970;
  assign n3972 = n3967 & n3968;
  assign n3973 = ~n3719 & n3966;
  assign n3974 = n3972 & n3973;
  assign po035 = ~n3971 | ~n3974;
  assign n3976 = n2677 & ~n2900;
  assign n3977 = ~n2902 & ~n3976;
  assign n3978 = pi029 & n1562;
  assign n3979 = n306 & n498;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = n329 & n480;
  assign n3982 = ~n3980 & n3981;
  assign n3983 = ~n360 & ~n3057;
  assign n3984 = ~n566 & n1504;
  assign n3985 = ~n2915 & ~n3226;
  assign n3986 = ~n3984 & n3985;
  assign n3987 = ~n3365 & n3986;
  assign n3988 = pi039 & n3542;
  assign n3989 = ~n3168 & ~n3988;
  assign n3990 = ~n2093 & n3989;
  assign n3991 = ~n3982 & n3990;
  assign n3992 = n3977 & n3991;
  assign n3993 = n3987 & n3992;
  assign n3994 = ~n3983 & n3993;
  assign n3995 = n638 & n1873;
  assign n3996 = n1073 & n3995;
  assign n3997 = ~n3629 & ~n3996;
  assign n3998 = n3649 & n3997;
  assign n3999 = n740 & n2684;
  assign n4000 = ~n528 & ~n2335;
  assign n4001 = ~n2001 & n4000;
  assign n4002 = ~pi001 & ~n4001;
  assign n4003 = ~n3999 & ~n4002;
  assign n4004 = ~pi007 & ~n4003;
  assign n4005 = ~n2993 & ~n3176;
  assign n4006 = n646 & n3037;
  assign n4007 = n2097 & n2961;
  assign n4008 = ~n722 & n2957;
  assign n4009 = n1172 & n1849;
  assign n4010 = pi013 & n3239;
  assign n4011 = pi012 & n1006;
  assign n4012 = n1749 & ~n4011;
  assign n4013 = n550 & n957;
  assign n4014 = ~n2263 & ~n4013;
  assign n4015 = n335 & ~n4014;
  assign n4016 = n2050 & n2600;
  assign n4017 = ~n2556 & ~n4016;
  assign n4018 = n299 & ~n4017;
  assign n4019 = ~n630 & ~n1076;
  assign n4020 = n3889 & ~n4019;
  assign n4021 = n320 & n3229;
  assign n4022 = ~pi029 & n533;
  assign n4023 = ~n532 & ~n4022;
  assign n4024 = ~n537 & ~n771;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = n733 & n2600;
  assign n4027 = n479 & n555;
  assign n4028 = n292 & n2025;
  assign n4029 = pi003 & n369;
  assign n4030 = n2000 & n4029;
  assign n4031 = n938 & n1490;
  assign n4032 = n1344 & n2619;
  assign n4033 = n1674 & ~n1746;
  assign n4034 = n944 & n4033;
  assign n4035 = n293 & ~n2941;
  assign n4036 = ~n2994 & ~n2996;
  assign n4037 = n1243 & n2798;
  assign n4038 = n4036 & ~n4037;
  assign n4039 = ~n4035 & n4038;
  assign n4040 = n345 & ~n4039;
  assign n4041 = ~pi021 & ~n3617;
  assign n4042 = n1873 & ~n4041;
  assign n4043 = ~n3622 & n4042;
  assign n4044 = n996 & ~n3172;
  assign n4045 = n1002 & n4044;
  assign n4046 = ~n990 & ~n4045;
  assign n4047 = pi013 & n2575;
  assign n4048 = pi029 & n4047;
  assign n4049 = ~n1242 & ~n1688;
  assign n4050 = n644 & ~n4049;
  assign n4051 = n3589 & ~n4050;
  assign n4052 = ~n3635 & n4051;
  assign n4053 = ~n3016 & n3269;
  assign n4054 = n4052 & ~n4053;
  assign n4055 = ~n3259 & n3593;
  assign n4056 = n4054 & n4055;
  assign n4057 = n1729 & n2575;
  assign n4058 = pi012 & n653;
  assign n4059 = n798 & n1699;
  assign n4060 = n4058 & n4059;
  assign n4061 = ~n734 & ~n1760;
  assign n4062 = pi014 & ~n4061;
  assign n4063 = n1465 & n3874;
  assign n4064 = n492 & ~n4063;
  assign n4065 = n1702 & n2623;
  assign n4066 = ~n2357 & ~n2367;
  assign n4067 = n329 & ~n4066;
  assign n4068 = ~pi088 & n293;
  assign n4069 = n521 & n4068;
  assign n4070 = ~n2589 & ~n4069;
  assign n4071 = ~n4067 & n4070;
  assign n4072 = ~n594 & ~n1528;
  assign n4073 = n677 & n692;
  assign n4074 = n771 & n1699;
  assign n4075 = n3473 & n4074;
  assign n4076 = ~n4073 & ~n4075;
  assign n4077 = ~pi015 & ~n4076;
  assign n4078 = n4072 & ~n4077;
  assign n4079 = n627 & n2029;
  assign n4080 = n332 & ~n584;
  assign n4081 = ~n680 & ~n4080;
  assign n4082 = n959 & ~n4081;
  assign n4083 = n1718 & n1780;
  assign n4084 = ~n3770 & ~n4083;
  assign n4085 = ~n4082 & n4084;
  assign n4086 = ~n3350 & n4085;
  assign n4087 = n960 & ~n4086;
  assign n4088 = ~n304 & ~n3312;
  assign n4089 = n854 & ~n4088;
  assign n4090 = ~pi013 & n3367;
  assign n4091 = ~n4087 & ~n4089;
  assign n4092 = ~n4090 & n4091;
  assign n4093 = n329 & ~n4092;
  assign n4094 = n290 & n2058;
  assign n4095 = ~n459 & ~n4094;
  assign n4096 = ~n2487 & n4095;
  assign n4097 = n451 & ~n4096;
  assign n4098 = ~n611 & ~n4079;
  assign n4099 = ~n4097 & n4098;
  assign n4100 = ~n4093 & n4099;
  assign n4101 = ~n2843 & n3840;
  assign n4102 = pi004 & ~n501;
  assign n4103 = n492 & n957;
  assign n4104 = ~n502 & n4103;
  assign n4105 = ~n4102 & n4104;
  assign n4106 = n427 & n511;
  assign n4107 = ~n1162 & ~n4106;
  assign n4108 = n576 & ~n4107;
  assign n4109 = n642 & n1870;
  assign n4110 = n1080 & n4109;
  assign n4111 = ~n4108 & ~n4110;
  assign n4112 = ~n1017 & n4111;
  assign n4113 = ~n4105 & n4112;
  assign n4114 = n2379 & n4113;
  assign n4115 = ~n2830 & n4114;
  assign n4116 = pi013 & ~n449;
  assign n4117 = n2531 & n4116;
  assign n4118 = ~pi010 & n3489;
  assign n4119 = n1011 & n2530;
  assign n4120 = ~n3678 & ~n4119;
  assign n4121 = ~n4117 & n4120;
  assign n4122 = ~n4118 & n4121;
  assign n4123 = ~n1325 & ~n1752;
  assign n4124 = n329 & n692;
  assign n4125 = n2182 & ~n4124;
  assign n4126 = n4123 & n4125;
  assign n4127 = n3295 & ~n4126;
  assign n4128 = n771 & n1724;
  assign n4129 = n1671 & n4128;
  assign n4130 = n643 & n778;
  assign n4131 = n338 & n405;
  assign n4132 = n376 & n2008;
  assign n4133 = n332 & n2114;
  assign n4134 = ~n4131 & ~n4132;
  assign n4135 = ~n2303 & n4134;
  assign n4136 = ~n4130 & n4135;
  assign n4137 = ~n4133 & n4136;
  assign n4138 = n369 & n550;
  assign n4139 = ~n762 & ~n4138;
  assign n4140 = n336 & ~n4139;
  assign n4141 = ~n567 & n1428;
  assign n4142 = n949 & n4141;
  assign n4143 = n1590 & n3642;
  assign n4144 = n2777 & n3840;
  assign n4145 = n630 & n4144;
  assign n4146 = ~n301 & ~n1704;
  assign n4147 = n304 & ~n4146;
  assign n4148 = ~pi006 & n689;
  assign n4149 = ~n3866 & ~n4148;
  assign n4150 = ~n1032 & n4149;
  assign n4151 = pi015 & ~n4150;
  assign n4152 = pi013 & n584;
  assign n4153 = n653 & ~n722;
  assign n4154 = ~n1033 & ~n4152;
  assign n4155 = ~n4153 & n4154;
  assign n4156 = n1753 & ~n4155;
  assign n4157 = n329 & n3301;
  assign n4158 = ~n2713 & ~n4157;
  assign n4159 = n1696 & ~n4158;
  assign n4160 = pi011 & n1987;
  assign n4161 = n791 & ~n3110;
  assign n4162 = n3730 & ~n4161;
  assign n4163 = n361 & ~n3087;
  assign n4164 = n1376 & n2388;
  assign n4165 = ~pi020 & n4164;
  assign n4166 = n606 & n2521;
  assign n4167 = ~n3472 & ~n4166;
  assign n4168 = n2831 & n2837;
  assign n4169 = pi065 & n2572;
  assign n4170 = ~n360 & n798;
  assign n4171 = n4169 & n4170;
  assign n4172 = n644 & n791;
  assign n4173 = n2571 & n4172;
  assign n4174 = ~n4171 & ~n4173;
  assign n4175 = n1376 & n2720;
  assign n4176 = n4174 & ~n4175;
  assign n4177 = ~n4168 & n4176;
  assign n4178 = n3837 & n4177;
  assign n4179 = ~n2582 & ~n3060;
  assign n4180 = ~n3539 & ~n3601;
  assign n4181 = n596 & n1590;
  assign n4182 = ~n3083 & ~n4181;
  assign n4183 = ~n382 & n4182;
  assign n4184 = n315 & ~n4183;
  assign n4185 = n4180 & ~n4184;
  assign n4186 = ~n1377 & n2880;
  assign n4187 = n4185 & ~n4186;
  assign n4188 = ~n1989 & ~n2029;
  assign n4189 = n1990 & ~n4188;
  assign n4190 = ~n1990 & ~n2522;
  assign n4191 = n1702 & ~n4190;
  assign n4192 = n853 & ~n3060;
  assign n4193 = n1228 & n2487;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = n1724 & ~n4194;
  assign n4196 = ~n4189 & ~n4195;
  assign n4197 = ~n4191 & n4196;
  assign n4198 = ~n2574 & n4197;
  assign n4199 = ~n4179 & n4198;
  assign n4200 = n4187 & n4199;
  assign n4201 = n3547 & n4200;
  assign n4202 = n1670 & n2911;
  assign n4203 = n898 & n4202;
  assign n4204 = n1671 & n2597;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = ~n1829 & n4205;
  assign n4207 = ~n468 & ~n3363;
  assign n4208 = n4206 & n4207;
  assign n4209 = n3373 & n4208;
  assign n4210 = n3708 & n4209;
  assign n4211 = n329 & ~n4210;
  assign n4212 = n825 & n993;
  assign n4213 = ~n2878 & ~n4212;
  assign n4214 = n514 & n646;
  assign n4215 = n417 & n4214;
  assign n4216 = n4213 & ~n4215;
  assign n4217 = n1071 & n3591;
  assign n4218 = n2772 & ~n2774;
  assign n4219 = n791 & ~n4218;
  assign n4220 = pi005 & n2331;
  assign n4221 = ~n2325 & ~n4220;
  assign n4222 = ~n474 & n3054;
  assign n4223 = ~n360 & n3061;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~n4219 & n4221;
  assign n4226 = n4224 & n4225;
  assign n4227 = n453 & n554;
  assign n4228 = ~n3215 & ~n4227;
  assign n4229 = ~pi004 & ~n4228;
  assign n4230 = pi009 & n625;
  assign n4231 = n2548 & n4230;
  assign n4232 = ~n4217 & ~n4229;
  assign n4233 = ~n4231 & n4232;
  assign n4234 = ~n2540 & n4233;
  assign n4235 = n4226 & n4234;
  assign n4236 = n714 & ~n1936;
  assign n4237 = ~n1294 & ~n1884;
  assign n4238 = n2677 & ~n4237;
  assign n4239 = n503 & n2792;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = ~n2710 & n4240;
  assign n4242 = ~n3746 & n4241;
  assign n4243 = n2767 & n4242;
  assign n4244 = ~n2661 & n2982;
  assign n4245 = n4243 & n4244;
  assign n4246 = ~n474 & n3045;
  assign n4247 = n1419 & n2234;
  assign n4248 = ~n569 & ~n2258;
  assign n4249 = n361 & ~n4248;
  assign n4250 = ~n972 & ~n1071;
  assign n4251 = n1975 & ~n4250;
  assign n4252 = n404 & n1922;
  assign n4253 = ~n3597 & ~n4252;
  assign n4254 = n551 & ~n4253;
  assign n4255 = ~n2288 & ~n4254;
  assign n4256 = ~n4251 & n4255;
  assign n4257 = n345 & n1387;
  assign n4258 = ~pi122 & n1049;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260 = n515 & ~n4259;
  assign n4261 = n492 & ~n2037;
  assign n4262 = ~n3100 & n4261;
  assign n4263 = ~n1435 & ~n2690;
  assign n4264 = n2663 & ~n4263;
  assign n4265 = n480 & n529;
  assign n4266 = ~n1398 & n4265;
  assign n4267 = n355 & n1404;
  assign n4268 = n668 & n1428;
  assign n4269 = n419 & n4268;
  assign n4270 = n353 & n1361;
  assign n4271 = n1399 & ~n4000;
  assign n4272 = ~pi122 & n2785;
  assign n4273 = ~n2800 & ~n4272;
  assign n4274 = ~n599 & n667;
  assign n4275 = n2234 & ~n4274;
  assign n4276 = ~n2230 & n4275;
  assign n4277 = ~n2298 & ~n4266;
  assign n4278 = n2328 & n4277;
  assign n4279 = ~n4269 & ~n4270;
  assign n4280 = ~n4271 & n4279;
  assign n4281 = ~n939 & n4278;
  assign n4282 = ~n4246 & n4281;
  assign n4283 = ~n4247 & n4280;
  assign n4284 = ~n4267 & n4283;
  assign n4285 = n1944 & n4282;
  assign n4286 = ~n3490 & ~n4236;
  assign n4287 = ~n4264 & ~n4276;
  assign n4288 = n4286 & n4287;
  assign n4289 = n4284 & n4285;
  assign n4290 = ~n3769 & n4256;
  assign n4291 = ~n4260 & ~n4262;
  assign n4292 = n4273 & n4291;
  assign n4293 = n4289 & n4290;
  assign n4294 = ~n4249 & n4288;
  assign n4295 = n4293 & n4294;
  assign n4296 = n4292 & n4295;
  assign n4297 = n4245 & n4296;
  assign n4298 = ~n4028 & ~n4030;
  assign n4299 = ~n4009 & n4298;
  assign n4300 = ~n4021 & ~n4025;
  assign n4301 = ~n4027 & n4300;
  assign n4302 = ~n1885 & n4299;
  assign n4303 = ~n3779 & ~n3842;
  assign n4304 = ~n4007 & ~n4008;
  assign n4305 = ~n4015 & ~n4026;
  assign n4306 = ~n4143 & ~n4159;
  assign n4307 = n4305 & n4306;
  assign n4308 = n4303 & n4304;
  assign n4309 = n4301 & n4302;
  assign n4310 = ~n1690 & ~n1973;
  assign n4311 = ~po123 & ~n3177;
  assign n4312 = ~n3614 & ~n4012;
  assign n4313 = ~n4018 & ~n4020;
  assign n4314 = ~n4032 & ~n4142;
  assign n4315 = ~n4160 & n4314;
  assign n4316 = n4312 & n4313;
  assign n4317 = n4310 & n4311;
  assign n4318 = n4308 & n4309;
  assign n4319 = ~n2598 & n4307;
  assign n4320 = n4005 & ~n4006;
  assign n4321 = ~n4031 & ~n4034;
  assign n4322 = ~n4127 & ~n4129;
  assign n4323 = n4137 & ~n4140;
  assign n4324 = ~n4151 & n4323;
  assign n4325 = n4321 & n4322;
  assign n4326 = n4319 & n4320;
  assign n4327 = n4317 & n4318;
  assign n4328 = n4315 & n4316;
  assign n4329 = n651 & n1721;
  assign n4330 = n3456 & n3612;
  assign n4331 = ~n3721 & ~n4004;
  assign n4332 = ~n4010 & ~n4060;
  assign n4333 = ~n4062 & ~n4147;
  assign n4334 = ~n4156 & ~n4165;
  assign n4335 = n4167 & n4334;
  assign n4336 = n4332 & n4333;
  assign n4337 = n4330 & n4331;
  assign n4338 = n4328 & n4329;
  assign n4339 = n4326 & n4327;
  assign n4340 = n4324 & n4325;
  assign n4341 = n691 & ~n4057;
  assign n4342 = ~n4065 & ~n4145;
  assign n4343 = n4341 & n4342;
  assign n4344 = n4339 & n4340;
  assign n4345 = n4337 & n4338;
  assign n4346 = n4335 & n4336;
  assign n4347 = n424 & ~n4048;
  assign n4348 = ~n4064 & ~n4101;
  assign n4349 = n4122 & ~n4163;
  assign n4350 = n4348 & n4349;
  assign n4351 = n4346 & n4347;
  assign n4352 = n4344 & n4345;
  assign n4353 = ~n2806 & n4343;
  assign n4354 = n2955 & n3799;
  assign n4355 = n3824 & n3998;
  assign n4356 = ~n4040 & ~n4043;
  assign n4357 = ~n4046 & n4071;
  assign n4358 = n4078 & n4100;
  assign n4359 = n4357 & n4358;
  assign n4360 = n4355 & n4356;
  assign n4361 = n4353 & n4354;
  assign n4362 = n4351 & n4352;
  assign n4363 = n3994 & n4350;
  assign n4364 = n4056 & n4115;
  assign n4365 = n4162 & n4364;
  assign n4366 = n4362 & n4363;
  assign n4367 = n4360 & n4361;
  assign n4368 = n3035 & n4359;
  assign n4369 = ~n4211 & n4368;
  assign n4370 = n4366 & n4367;
  assign n4371 = n4178 & n4365;
  assign n4372 = n4216 & n4235;
  assign n4373 = n4371 & n4372;
  assign n4374 = n4369 & n4370;
  assign n4375 = n4201 & n4297;
  assign n4376 = n4374 & n4375;
  assign n4377 = n4373 & n4376;
  assign po036 = ~n3162 | ~n4377;
  assign n4379 = n494 & n2702;
  assign n4380 = n2824 & ~n4379;
  assign n4381 = ~n1968 & n4380;
  assign n4382 = n1983 & n4381;
  assign n4383 = n1266 & ~n1285;
  assign n4384 = n1846 & n4383;
  assign n4385 = ~pi045 & pi122;
  assign n4386 = n1164 & n4385;
  assign n4387 = pi056 & n1136;
  assign n4388 = n4385 & ~n4387;
  assign n4389 = ~n811 & ~n4388;
  assign n4390 = ~n2861 & ~n4389;
  assign n4391 = ~n1166 & n1183;
  assign n4392 = ~n2105 & n4391;
  assign n4393 = ~pi045 & ~n4392;
  assign n4394 = n1147 & ~n1331;
  assign n4395 = ~n1193 & ~n4394;
  assign n4396 = n293 & n811;
  assign n4397 = ~n4395 & n4396;
  assign n4398 = n1205 & n1892;
  assign n4399 = ~pi056 & n306;
  assign n4400 = n4398 & n4399;
  assign n4401 = ~n4390 & ~n4400;
  assign n4402 = ~n4397 & n4401;
  assign n4403 = ~n4393 & n4402;
  assign n4404 = ~n4386 & n4403;
  assign n4405 = ~pi045 & n293;
  assign n4406 = pi022 & n4405;
  assign n4407 = n3068 & n4406;
  assign n4408 = n4404 & ~n4407;
  assign n4409 = pi006 & n1207;
  assign n4410 = n2866 & ~n4409;
  assign n4411 = ~pi045 & ~n4410;
  assign n4412 = n798 & ~n1229;
  assign n4413 = ~n4389 & n4412;
  assign n4414 = ~n4411 & ~n4413;
  assign n4415 = n332 & n439;
  assign n4416 = ~n584 & n4415;
  assign n4417 = n492 & ~n2102;
  assign n4418 = n1151 & ~n2860;
  assign n4419 = ~n1194 & n4418;
  assign n4420 = ~n1186 & n4419;
  assign n4421 = ~n1998 & n4420;
  assign n4422 = ~n2854 & n4421;
  assign n4423 = ~n4417 & n4422;
  assign n4424 = n4388 & ~n4423;
  assign n4425 = n744 & n993;
  assign n4426 = ~n1328 & ~n4425;
  assign n4427 = ~pi029 & n2646;
  assign n4428 = ~n4426 & n4427;
  assign n4429 = ~n4424 & ~n4428;
  assign n4430 = n1219 & n1228;
  assign n4431 = ~n1227 & ~n4430;
  assign n4432 = n2095 & n4431;
  assign n4433 = n3339 & n4432;
  assign n4434 = n363 & n575;
  assign n4435 = n460 & n673;
  assign n4436 = ~n799 & n1583;
  assign n4437 = pi022 & n3000;
  assign n4438 = n3235 & ~n4434;
  assign n4439 = ~n4436 & n4438;
  assign n4440 = ~n4437 & n4439;
  assign n4441 = n3795 & ~n4416;
  assign n4442 = ~n4435 & n4441;
  assign n4443 = n4440 & n4442;
  assign n4444 = n4414 & n4443;
  assign n4445 = n4433 & n4444;
  assign n4446 = n4408 & n4445;
  assign n4447 = n4429 & n4446;
  assign n4448 = n330 & n1441;
  assign n4449 = n1294 & n1306;
  assign n4450 = n1437 & n4449;
  assign n4451 = n302 & n823;
  assign n4452 = ~n1437 & n2590;
  assign n4453 = ~n332 & n3894;
  assign n4454 = ~n750 & n802;
  assign n4455 = ~pi028 & ~pi108;
  assign n4456 = n4454 & ~n4455;
  assign n4457 = ~pi019 & n1421;
  assign n4458 = ~pi074 & n3890;
  assign n4459 = n1008 & n1775;
  assign n4460 = n568 & n1975;
  assign n4461 = n798 & n1436;
  assign n4462 = n1884 & ~n2614;
  assign n4463 = ~pi023 & n1520;
  assign n4464 = ~n1887 & ~n4462;
  assign n4465 = ~n4461 & ~n4463;
  assign n4466 = n4464 & n4465;
  assign n4467 = ~n590 & ~n2961;
  assign n4468 = n336 & ~n4467;
  assign n4469 = ~n568 & ~n2411;
  assign n4470 = n429 & ~n4469;
  assign n4471 = ~n341 & ~n823;
  assign n4472 = pi015 & ~n4471;
  assign n4473 = pi012 & n467;
  assign n4474 = ~n1775 & n4473;
  assign n4475 = ~n1468 & ~n3869;
  assign n4476 = n1376 & ~n4475;
  assign n4477 = n1376 & n1464;
  assign n4478 = ~n649 & ~n4477;
  assign n4479 = ~n710 & ~n2957;
  assign n4480 = n493 & ~n4479;
  assign n4481 = n332 & n726;
  assign n4482 = n729 & ~n4481;
  assign n4483 = ~pi015 & ~n4482;
  assign n4484 = n1428 & n2256;
  assign n4485 = pi007 & ~pi108;
  assign n4486 = n749 & n4485;
  assign n4487 = ~n1623 & ~n4486;
  assign n4488 = ~n807 & n4487;
  assign n4489 = ~n4484 & n4488;
  assign n4490 = n492 & ~n4489;
  assign n4491 = ~n1474 & ~n1591;
  assign n4492 = n492 & n577;
  assign n4493 = ~n2110 & ~n4492;
  assign n4494 = n2411 & ~n4493;
  assign n4495 = ~n1336 & ~n1916;
  assign n4496 = ~n470 & n4495;
  assign n4497 = ~n3109 & n4496;
  assign n4498 = n330 & ~n4497;
  assign n4499 = ~n446 & ~n497;
  assign n4500 = ~n641 & ~n2318;
  assign n4501 = ~n4448 & ~n4451;
  assign n4502 = ~n4452 & ~n4470;
  assign n4503 = n4501 & n4502;
  assign n4504 = n4499 & n4500;
  assign n4505 = ~n4450 & ~n4459;
  assign n4506 = ~n4468 & n4505;
  assign n4507 = n4503 & n4504;
  assign n4508 = ~n365 & ~n3906;
  assign n4509 = ~n4453 & ~n4456;
  assign n4510 = ~n4458 & ~n4472;
  assign n4511 = n4509 & n4510;
  assign n4512 = n4507 & n4508;
  assign n4513 = ~n4460 & n4506;
  assign n4514 = ~n4474 & ~n4480;
  assign n4515 = ~n4483 & ~n4494;
  assign n4516 = n4514 & n4515;
  assign n4517 = n4512 & n4513;
  assign n4518 = n3287 & n4511;
  assign n4519 = n3742 & ~n4457;
  assign n4520 = ~n4476 & n4478;
  assign n4521 = ~n4490 & n4520;
  assign n4522 = n4518 & n4519;
  assign n4523 = n4516 & n4517;
  assign n4524 = n3767 & n4466;
  assign n4525 = n4523 & n4524;
  assign n4526 = n4521 & n4522;
  assign n4527 = ~n942 & ~n2261;
  assign n4528 = n4491 & n4527;
  assign n4529 = n4525 & n4526;
  assign n4530 = n858 & n1341;
  assign n4531 = n4529 & n4530;
  assign n4532 = n4384 & n4528;
  assign n4533 = ~n4498 & n4532;
  assign n4534 = n4531 & n4533;
  assign n4535 = n4447 & n4534;
  assign po037 = ~n4382 | ~n4535;
  assign n4537 = ~n1030 & ~n1228;
  assign n4538 = n2035 & ~n4537;
  assign n4539 = n1338 & ~n3528;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = n1320 & n4540;
  assign n4542 = n2542 & n4541;
  assign n4543 = ~n2370 & n4542;
  assign n4544 = ~n790 & n3110;
  assign n4545 = n4496 & n4544;
  assign n4546 = n330 & ~n4545;
  assign n4547 = n704 & n1772;
  assign n4548 = ~n1744 & ~n3295;
  assign n4549 = n1011 & ~n4548;
  assign n4550 = n493 & n2097;
  assign n4551 = n444 & n4550;
  assign n4552 = pi013 & n823;
  assign n4553 = ~n520 & ~n2505;
  assign n4554 = n518 & ~n4553;
  assign n4555 = n302 & n340;
  assign n4556 = n315 & n2008;
  assign n4557 = ~pi074 & n4020;
  assign n4558 = n368 & ~n2113;
  assign n4559 = ~pi023 & n567;
  assign n4560 = n315 & n636;
  assign n4561 = ~n4559 & n4560;
  assign n4562 = n1295 & n4561;
  assign n4563 = pi015 & n442;
  assign n4564 = n723 & n4563;
  assign n4565 = n521 & n957;
  assign n4566 = n957 & n2005;
  assign n4567 = pi014 & ~n332;
  assign n4568 = ~n727 & n4567;
  assign n4569 = n733 & n4568;
  assign n4570 = ~pi002 & ~n1922;
  assign n4571 = ~pi005 & ~n4570;
  assign n4572 = ~n308 & ~n4571;
  assign n4573 = n554 & ~n4572;
  assign n4574 = n411 & n2415;
  assign n4575 = n348 & n1712;
  assign n4576 = n369 & ~n2265;
  assign n4577 = n607 & n902;
  assign n4578 = n2548 & n4577;
  assign n4579 = n506 & n1076;
  assign n4580 = pi012 & n1416;
  assign n4581 = n1715 & n4181;
  assign n4582 = pi022 & n1388;
  assign n4583 = n638 & n773;
  assign n4584 = ~n2961 & ~n4583;
  assign n4585 = ~n4582 & n4584;
  assign n4586 = n315 & ~n4585;
  assign n4587 = n598 & n2528;
  assign n4588 = ~n4457 & ~n4587;
  assign n4589 = ~n3759 & n4588;
  assign n4590 = ~n1388 & n2259;
  assign n4591 = n361 & ~n4590;
  assign n4592 = ~pi022 & n668;
  assign n4593 = n698 & n4592;
  assign n4594 = n938 & ~n2267;
  assign n4595 = n293 & n965;
  assign n4596 = n319 & n4595;
  assign n4597 = ~n3206 & ~n4596;
  assign n4598 = ~n4594 & n4597;
  assign n4599 = ~n4593 & n4598;
  assign n4600 = ~n2194 & n4599;
  assign n4601 = ~n1286 & ~n1541;
  assign n4602 = ~n3289 & n4601;
  assign n4603 = pi015 & n3679;
  assign n4604 = ~n303 & n2532;
  assign n4605 = ~pi018 & n1766;
  assign n4606 = ~n1386 & ~n4605;
  assign n4607 = ~pi023 & ~n4606;
  assign n4608 = n1069 & n1392;
  assign n4609 = n410 & n1275;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = n1385 & ~n4610;
  assign n4612 = ~n299 & ~n1673;
  assign n4613 = n1697 & ~n4612;
  assign n4614 = ~n2522 & ~n4613;
  assign n4615 = n852 & ~n4614;
  assign n4616 = pi018 & n1765;
  assign n4617 = ~n2659 & ~n4448;
  assign n4618 = ~n303 & n708;
  assign n4619 = ~n681 & ~n3229;
  assign n4620 = n1749 & ~n4619;
  assign n4621 = ~pi021 & n3624;
  assign n4622 = ~n1876 & ~n4621;
  assign n4623 = ~n2078 & n4622;
  assign n4624 = ~pi018 & ~n4623;
  assign n4625 = ~n1901 & ~n2244;
  assign n4626 = n2248 & n4625;
  assign n4627 = ~n360 & ~n4626;
  assign n4628 = ~n2227 & ~n2229;
  assign n4629 = n2234 & ~n4628;
  assign n4630 = n858 & ~n1727;
  assign n4631 = pi023 & n2471;
  assign n4632 = n1752 & n4202;
  assign n4633 = ~n448 & n1659;
  assign n4634 = n1673 & n4633;
  assign n4635 = ~n3454 & ~n4634;
  assign n4636 = ~pi012 & ~n4635;
  assign n4637 = ~n2554 & ~n4632;
  assign n4638 = ~n4636 & n4637;
  assign n4639 = ~pi015 & ~n4638;
  assign n4640 = n466 & n2600;
  assign n4641 = n678 & n1033;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~n4164 & n4642;
  assign n4644 = ~n2508 & ~n4556;
  assign n4645 = ~n634 & n4644;
  assign n4646 = ~n690 & ~n1572;
  assign n4647 = ~n1883 & ~n1931;
  assign n4648 = ~n4565 & ~n4573;
  assign n4649 = n4647 & n4648;
  assign n4650 = n4645 & n4646;
  assign n4651 = ~n728 & ~n2266;
  assign n4652 = ~n3176 & ~n4551;
  assign n4653 = ~n4552 & ~n4554;
  assign n4654 = ~n4555 & ~n4562;
  assign n4655 = ~n4564 & ~n4566;
  assign n4656 = ~n4569 & ~n4576;
  assign n4657 = n4655 & n4656;
  assign n4658 = n4653 & n4654;
  assign n4659 = n4651 & n4652;
  assign n4660 = n4649 & n4650;
  assign n4661 = ~n504 & ~n4454;
  assign n4662 = ~n4558 & ~n4574;
  assign n4663 = ~n4578 & ~n4580;
  assign n4664 = ~n4581 & ~n4620;
  assign n4665 = n4663 & n4664;
  assign n4666 = n4661 & n4662;
  assign n4667 = n4659 & n4660;
  assign n4668 = n4657 & n4658;
  assign n4669 = ~n409 & n650;
  assign n4670 = ~n951 & n2591;
  assign n4671 = ~n2594 & ~n2602;
  assign n4672 = ~n3481 & ~n4119;
  assign n4673 = n4137 & ~n4547;
  assign n4674 = ~n4557 & ~n4575;
  assign n4675 = ~n4579 & ~n4618;
  assign n4676 = n4674 & n4675;
  assign n4677 = n4672 & n4673;
  assign n4678 = n4670 & n4671;
  assign n4679 = n4668 & n4669;
  assign n4680 = n4666 & n4667;
  assign n4681 = ~n2358 & n4665;
  assign n4682 = n2599 & ~n4549;
  assign n4683 = ~n4603 & ~n4616;
  assign n4684 = ~n4629 & n4643;
  assign n4685 = n4683 & n4684;
  assign n4686 = n4681 & n4682;
  assign n4687 = n4679 & n4680;
  assign n4688 = n4677 & n4678;
  assign n4689 = n613 & n4676;
  assign n4690 = n701 & ~n1395;
  assign n4691 = n1762 & n1888;
  assign n4692 = ~n1980 & n4256;
  assign n4693 = ~n4604 & ~n4607;
  assign n4694 = ~n4611 & n4617;
  assign n4695 = n4693 & n4694;
  assign n4696 = n4691 & n4692;
  assign n4697 = n4689 & n4690;
  assign n4698 = n4687 & n4688;
  assign n4699 = n4685 & n4686;
  assign n4700 = n872 & ~n4586;
  assign n4701 = n4600 & ~n4615;
  assign n4702 = ~n4631 & n4701;
  assign n4703 = n4699 & n4700;
  assign n4704 = n4697 & n4698;
  assign n4705 = n4695 & n4696;
  assign n4706 = n367 & n4589;
  assign n4707 = ~n4591 & n4602;
  assign n4708 = ~n4624 & ~n4639;
  assign n4709 = n4707 & n4708;
  assign n4710 = n4705 & n4706;
  assign n4711 = n4703 & n4704;
  assign n4712 = n946 & n4702;
  assign n4713 = n2354 & ~n2468;
  assign n4714 = ~n3292 & n4713;
  assign n4715 = n4711 & n4712;
  assign n4716 = n4709 & n4710;
  assign n4717 = n1864 & ~n4546;
  assign n4718 = ~n4627 & n4630;
  assign n4719 = n4717 & n4718;
  assign n4720 = n4715 & n4716;
  assign n4721 = n4714 & n4720;
  assign n4722 = n3386 & n4719;
  assign n4723 = n4721 & n4722;
  assign n4724 = n4447 & n4723;
  assign n4725 = n4543 & n4724;
  assign po038 = ~n4381 | ~n4725;
  assign n4727 = n476 & n938;
  assign n4728 = n408 & n1501;
  assign n4729 = n2592 & ~n4728;
  assign n4730 = ~pi029 & n1502;
  assign n4731 = ~n1311 & ~n3999;
  assign n4732 = n778 & n1074;
  assign n4733 = n555 & ~n2965;
  assign n4734 = ~n2508 & ~n4727;
  assign n4735 = ~n4733 & n4734;
  assign n4736 = ~n4449 & n4735;
  assign n4737 = ~n4732 & n4736;
  assign n4738 = ~n557 & n4737;
  assign n4739 = n1273 & n4731;
  assign n4740 = n4738 & n4739;
  assign n4741 = n4729 & n4740;
  assign n4742 = ~n4730 & n4741;
  assign po039 = ~n4466 | ~n4742;
  assign n4744 = n402 & n791;
  assign n4745 = ~n360 & n3056;
  assign n4746 = n1463 & ~n2908;
  assign n4747 = ~n571 & n604;
  assign n4748 = n604 & n1886;
  assign n4749 = ~n740 & ~n1093;
  assign n4750 = ~n330 & n1346;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = n1345 & n4751;
  assign n4753 = ~n4748 & ~n4752;
  assign n4754 = ~n798 & ~n802;
  assign n4755 = n1583 & ~n4754;
  assign n4756 = n4005 & ~n4755;
  assign n4757 = ~n4746 & n4756;
  assign n4758 = ~n2909 & ~n4747;
  assign n4759 = n4757 & n4758;
  assign n4760 = n4753 & n4759;
  assign n4761 = ~n4745 & n4760;
  assign n4762 = ~n3033 & n4761;
  assign n4763 = n3118 & ~n3292;
  assign n4764 = n4762 & n4763;
  assign n4765 = n2684 & ~n3733;
  assign n4766 = ~n2771 & ~n2774;
  assign n4767 = n791 & ~n4766;
  assign n4768 = n3103 & n3814;
  assign n4769 = n416 & ~n990;
  assign n4770 = n570 & n4769;
  assign n4771 = n329 & n3278;
  assign n4772 = n450 & n492;
  assign n4773 = n459 & n4772;
  assign n4774 = ~n3184 & ~n4771;
  assign n4775 = ~n4773 & n4774;
  assign n4776 = n1847 & n1849;
  assign n4777 = n416 & n477;
  assign n4778 = ~n997 & ~n4777;
  assign n4779 = n330 & ~n4778;
  assign n4780 = ~n2873 & ~n4776;
  assign n4781 = ~n1269 & n4780;
  assign n4782 = ~n4744 & ~n4765;
  assign n4783 = n4781 & n4782;
  assign n4784 = ~n4770 & ~n4779;
  assign n4785 = n4783 & n4784;
  assign n4786 = n4775 & n4785;
  assign n4787 = ~n3728 & ~n4767;
  assign n4788 = ~n4768 & n4787;
  assign n4789 = n1890 & n4786;
  assign n4790 = n4788 & n4789;
  assign n4791 = n1340 & n1947;
  assign n4792 = n4790 & n4791;
  assign n4793 = n2240 & n4792;
  assign n4794 = n4178 & n4764;
  assign n4795 = n4793 & n4794;
  assign n4796 = n1093 & n1699;
  assign n4797 = n1730 & n4796;
  assign n4798 = n510 & ~n667;
  assign n4799 = n1685 & n4798;
  assign n4800 = ~n1690 & ~n4799;
  assign n4801 = ~n1876 & n4800;
  assign n4802 = n3998 & n4801;
  assign n4803 = n4056 & n4802;
  assign n4804 = ~n1916 & n3708;
  assign n4805 = ~n2357 & ~n3300;
  assign n4806 = n4804 & n4805;
  assign n4807 = n329 & ~n4806;
  assign n4808 = ~n790 & ~n2774;
  assign n4809 = n4045 & n4808;
  assign n4810 = n330 & ~n4809;
  assign n4811 = ~pi013 & n2575;
  assign n4812 = ~n3771 & ~n4083;
  assign n4813 = ~n3772 & n4812;
  assign n4814 = n1786 & ~n4813;
  assign n4815 = ~n4811 & ~n4814;
  assign n4816 = ~pi029 & ~n4815;
  assign n4817 = ~n2988 & ~n2996;
  assign n4818 = n345 & ~n4817;
  assign n4819 = pi029 & ~n464;
  assign n4820 = ~pi029 & ~n1033;
  assign n4821 = ~n2029 & n4820;
  assign n4822 = ~n4819 & ~n4821;
  assign n4823 = ~n1724 & ~n4822;
  assign n4824 = n1753 & ~n4823;
  assign n4825 = n3278 & n4170;
  assign n4826 = n529 & ~n2931;
  assign n4827 = pi001 & n1385;
  assign n4828 = ~n4826 & ~n4827;
  assign n4829 = n1396 & ~n4828;
  assign n4830 = n1696 & n4157;
  assign n4831 = ~n1693 & ~n1704;
  assign n4832 = n304 & ~n4831;
  assign n4833 = n1699 & ~n3060;
  assign n4834 = n3473 & n4833;
  assign n4835 = n2903 & n4080;
  assign n4836 = ~n4272 & ~n4835;
  assign n4837 = ~n2008 & ~n2057;
  assign n4838 = ~n1719 & ~n4632;
  assign n4839 = n2599 & ~n4018;
  assign n4840 = ~n1749 & n4839;
  assign n4841 = n4122 & n4840;
  assign n4842 = pi013 & n4079;
  assign n4843 = ~n703 & ~n1525;
  assign n4844 = n1704 & ~n4843;
  assign n4845 = ~n3532 & ~n4844;
  assign n4846 = ~pi014 & ~n4845;
  assign n4847 = n329 & n3353;
  assign n4848 = n854 & n1668;
  assign n4849 = ~n2689 & ~n4263;
  assign n4850 = ~n3473 & ~n4128;
  assign n4851 = n1671 & ~n4850;
  assign n4852 = n2388 & ~n2908;
  assign n4853 = ~n2521 & ~n2550;
  assign n4854 = n606 & ~n4853;
  assign n4855 = ~n1987 & ~n4854;
  assign n4856 = n3525 & n4855;
  assign n4857 = ~n4852 & n4856;
  assign n4858 = n780 & ~n781;
  assign n4859 = n471 & n4858;
  assign n4860 = ~n1829 & ~n3367;
  assign n4861 = ~n2367 & n4860;
  assign n4862 = n3373 & n4861;
  assign n4863 = n4859 & n4862;
  assign n4864 = n492 & ~n4863;
  assign n4865 = n3463 & ~n4110;
  assign n4866 = ~n4829 & ~n4830;
  assign n4867 = n4865 & n4866;
  assign n4868 = n3486 & ~n4825;
  assign n4869 = n4867 & n4868;
  assign n4870 = n4838 & ~n4842;
  assign n4871 = ~n4847 & ~n4848;
  assign n4872 = ~n4851 & n4871;
  assign n4873 = n4869 & n4870;
  assign n4874 = n2322 & n2377;
  assign n4875 = ~n4797 & ~n4824;
  assign n4876 = ~n4834 & n4837;
  assign n4877 = ~n4849 & n4876;
  assign n4878 = n4874 & n4875;
  assign n4879 = n4872 & n4873;
  assign n4880 = ~n1327 & n2312;
  assign n4881 = ~n4818 & ~n4832;
  assign n4882 = n4836 & ~n4846;
  assign n4883 = n4881 & n4882;
  assign n4884 = n4879 & n4880;
  assign n4885 = n4877 & n4878;
  assign n4886 = ~n1508 & ~n1756;
  assign n4887 = ~n1792 & ~n2235;
  assign n4888 = n4886 & n4887;
  assign n4889 = n4884 & n4885;
  assign n4890 = ~n4816 & n4883;
  assign n4891 = n4841 & n4890;
  assign n4892 = n4888 & n4889;
  assign n4893 = n2807 & n3626;
  assign n4894 = n4224 & ~n4810;
  assign n4895 = n4857 & n4894;
  assign n4896 = n4892 & n4893;
  assign n4897 = n4803 & n4891;
  assign n4898 = ~n4864 & n4897;
  assign n4899 = n4895 & n4896;
  assign n4900 = n4245 & ~n4807;
  assign n4901 = n4899 & n4900;
  assign n4902 = n4201 & n4898;
  assign n4903 = n4901 & n4902;
  assign n4904 = n4795 & n4903;
  assign po040 = ~n4543 | ~n4904;
  assign n4906 = n329 & ~n4804;
  assign n4907 = n442 & n1754;
  assign n4908 = ~n1033 & ~n1940;
  assign n4909 = n2623 & ~n4908;
  assign n4910 = ~n1724 & ~n1729;
  assign n4911 = n854 & ~n4910;
  assign n4912 = n303 & ~n722;
  assign n4913 = n3347 & n4912;
  assign n4914 = ~n4911 & ~n4913;
  assign n4915 = n492 & ~n4914;
  assign n4916 = ~pi029 & n360;
  assign n4917 = ~n2804 & ~n4916;
  assign n4918 = n439 & n450;
  assign n4919 = ~n3259 & ~n3638;
  assign n4920 = ~n3043 & ~n4825;
  assign n4921 = ~n1520 & ~n4849;
  assign n4922 = ~n2487 & ~n4094;
  assign n4923 = n3331 & ~n4922;
  assign n4924 = ~n3772 & n4086;
  assign n4925 = n1787 & ~n4924;
  assign n4926 = n532 & n1093;
  assign n4927 = pi029 & ~n2779;
  assign n4928 = n3547 & ~n4927;
  assign n4929 = ~n533 & n4809;
  assign n4930 = n330 & ~n4929;
  assign n4931 = n1664 & ~n2578;
  assign n4932 = ~n2388 & n4859;
  assign n4933 = ~n2357 & n4861;
  assign n4934 = n4931 & n4933;
  assign n4935 = n4932 & n4934;
  assign n4936 = n492 & ~n4935;
  assign n4937 = ~n2705 & ~n4926;
  assign n4938 = ~n3524 & n4937;
  assign n4939 = ~n4918 & ~n4923;
  assign n4940 = n4938 & n4939;
  assign n4941 = ~n2881 & ~n2971;
  assign n4942 = n3863 & ~n4925;
  assign n4943 = n4941 & n4942;
  assign n4944 = ~n4907 & n4940;
  assign n4945 = ~n4909 & ~n4915;
  assign n4946 = n4919 & n4921;
  assign n4947 = n4945 & n4946;
  assign n4948 = n4943 & n4944;
  assign n4949 = ~n4917 & n4920;
  assign n4950 = n4948 & n4949;
  assign n4951 = ~n4223 & n4947;
  assign n4952 = n4950 & n4951;
  assign n4953 = n4243 & n4952;
  assign n4954 = ~n4906 & ~n4930;
  assign n4955 = ~n4936 & n4954;
  assign n4956 = n4928 & n4953;
  assign n4957 = n4955 & n4956;
  assign n4958 = n3015 & n4957;
  assign n4959 = n4542 & n4795;
  assign po041 = ~n4958 | ~n4959;
  assign n4961 = n682 & n1834;
  assign n4962 = ~pi012 & ~n448;
  assign n4963 = n665 & n4962;
  assign n4964 = n1696 & n2704;
  assign n4965 = ~n3382 & ~n4964;
  assign n4966 = ~n4963 & n4965;
  assign n4967 = n3157 & n4966;
  assign n4968 = ~n3285 & ~n4961;
  assign n4969 = n1046 & n4968;
  assign n4970 = n4967 & n4969;
  assign n4971 = ~n1511 & ~n2714;
  assign n4972 = n2064 & n4971;
  assign n4973 = n3288 & n4972;
  assign n4974 = n4970 & n4973;
  assign n4975 = n3362 & n4974;
  assign n4976 = n1718 & n1754;
  assign n4977 = ~n2834 & n4144;
  assign n4978 = n798 & n1029;
  assign n4979 = ~n2881 & ~n4976;
  assign n4980 = ~n4977 & ~n4978;
  assign n4981 = n4979 & n4980;
  assign n4982 = ~pi060 & n2661;
  assign n4983 = n652 & n1024;
  assign n4984 = pi069 & n4983;
  assign n4985 = ~n4982 & ~n4984;
  assign n4986 = n460 & n1668;
  assign n4987 = n740 & ~n4045;
  assign n4988 = ~pi013 & n4079;
  assign n4989 = ~n440 & ~n4988;
  assign n4990 = n345 & n2988;
  assign n4991 = n2802 & ~n4990;
  assign n4992 = n961 & n4080;
  assign n4993 = n1912 & ~n4992;
  assign n4994 = n330 & ~n4993;
  assign n4995 = ~n2597 & ~n4124;
  assign n4996 = n3295 & ~n4995;
  assign n4997 = ~n1375 & ~n1517;
  assign n4998 = n2669 & ~n4997;
  assign n4999 = n345 & n2243;
  assign n5000 = n1092 & n2692;
  assign n5001 = pi027 & n5000;
  assign n5002 = n703 & n2903;
  assign n5003 = ~n1025 & ~n5002;
  assign n5004 = pi012 & ~n5003;
  assign n5005 = n1223 & ~n1999;
  assign n5006 = n1233 & ~n2103;
  assign n5007 = n5005 & n5006;
  assign n5008 = n752 & n1455;
  assign n5009 = ~n4164 & ~n5008;
  assign n5010 = n798 & ~n4858;
  assign n5011 = n5009 & ~n5010;
  assign n5012 = n554 & ~n2067;
  assign n5013 = ~pi002 & n5012;
  assign n5014 = pi044 & pi122;
  assign n5015 = ~pi000 & ~n5014;
  assign n5016 = ~n4388 & ~n5015;
  assign n5017 = pi002 & n295;
  assign n5018 = n827 & n5017;
  assign n5019 = ~n5016 & n5018;
  assign n5020 = n2840 & n3840;
  assign n5021 = ~n1011 & ~n1325;
  assign n5022 = n439 & ~n5021;
  assign n5023 = n492 & ~n750;
  assign n5024 = n625 & n627;
  assign n5025 = ~n3899 & ~n4034;
  assign n5026 = n678 & n1718;
  assign n5027 = n442 & n621;
  assign n5028 = ~n2055 & n5027;
  assign n5029 = ~n5026 & ~n5028;
  assign n5030 = n2245 & ~n2785;
  assign n5031 = ~pi122 & ~n5030;
  assign n5032 = n1786 & ~n4812;
  assign n5033 = n1693 & n3312;
  assign n5034 = ~n1329 & ~n3999;
  assign n5035 = ~n5032 & n5034;
  assign n5036 = ~n3856 & ~n5033;
  assign n5037 = n5035 & n5036;
  assign n5038 = ~n2484 & ~n4067;
  assign n5039 = n433 & n5038;
  assign n5040 = n4803 & n5039;
  assign n5041 = ~n3363 & n3540;
  assign n5042 = n329 & ~n5041;
  assign n5043 = n3086 & n3091;
  assign n5044 = n2260 & n5043;
  assign n5045 = ~n3080 & n5044;
  assign n5046 = n361 & ~n5045;
  assign n5047 = ~n1092 & ~n2539;
  assign n5048 = n1228 & ~n5047;
  assign n5049 = n506 & n933;
  assign n5050 = n615 & n1071;
  assign n5051 = pi013 & n1416;
  assign n5052 = n339 & ~n1795;
  assign n5053 = ~n957 & ~n4068;
  assign n5054 = n521 & ~n5053;
  assign n5055 = n311 & n829;
  assign n5056 = pi013 & pi015;
  assign n5057 = ~n1007 & ~n5056;
  assign n5058 = pi006 & ~n5057;
  assign n5059 = n726 & n5058;
  assign n5060 = ~n966 & ~n2112;
  assign n5061 = n368 & ~n5060;
  assign n5062 = ~n3012 & ~n5052;
  assign n5063 = ~n5054 & ~n5055;
  assign n5064 = n5062 & n5063;
  assign n5065 = ~n446 & ~n5059;
  assign n5066 = n5064 & n5065;
  assign n5067 = ~n5051 & ~n5061;
  assign n5068 = n5066 & n5067;
  assign n5069 = ~n3892 & ~n4746;
  assign n5070 = ~n5049 & ~n5050;
  assign n5071 = n5069 & n5070;
  assign n5072 = ~n1421 & n5068;
  assign n5073 = n5071 & n5072;
  assign n5074 = ~n2278 & n5073;
  assign n5075 = n4600 & ~n5048;
  assign n5076 = n5074 & n5075;
  assign n5077 = ~n3007 & n5076;
  assign n5078 = ~n5046 & n5077;
  assign n5079 = n4541 & n5078;
  assign n5080 = ~n1153 & ~n1175;
  assign n5081 = n4419 & n5080;
  assign n5082 = n4388 & ~n5081;
  assign n5083 = ~n1087 & n3155;
  assign n5084 = ~pi029 & n797;
  assign n5085 = n801 & n5084;
  assign n5086 = pi028 & n5085;
  assign n5087 = n5083 & ~n5086;
  assign n5088 = n1328 & n4427;
  assign n5089 = ~n4411 & ~n5088;
  assign n5090 = n4408 & n5089;
  assign n5091 = ~n5013 & ~n5019;
  assign n5092 = ~n795 & n5091;
  assign n5093 = ~n1272 & n5092;
  assign n5094 = n2757 & ~n3727;
  assign n5095 = ~n4238 & ~n5020;
  assign n5096 = ~n5023 & ~n5024;
  assign n5097 = n5095 & n5096;
  assign n5098 = n5093 & n5094;
  assign n5099 = ~n4996 & ~n4999;
  assign n5100 = ~n5022 & n5099;
  assign n5101 = n5097 & n5098;
  assign n5102 = ~n857 & n1042;
  assign n5103 = ~n4461 & ~n4986;
  assign n5104 = n4989 & ~n4998;
  assign n5105 = n5025 & n5029;
  assign n5106 = n5104 & n5105;
  assign n5107 = n5102 & n5103;
  assign n5108 = n5100 & n5101;
  assign n5109 = n343 & n3341;
  assign n5110 = n3722 & n4753;
  assign n5111 = ~n4767 & n5110;
  assign n5112 = n5108 & n5109;
  assign n5113 = n5106 & n5107;
  assign n5114 = n614 & n2316;
  assign n5115 = ~n3041 & n4176;
  assign n5116 = ~n4184 & n4985;
  assign n5117 = n4991 & ~n5001;
  assign n5118 = ~n5004 & ~n5031;
  assign n5119 = n5037 & n5118;
  assign n5120 = n5116 & n5117;
  assign n5121 = n5114 & n5115;
  assign n5122 = n5112 & n5113;
  assign n5123 = n3052 & n5111;
  assign n5124 = n4114 & n4981;
  assign n5125 = ~n4987 & ~n4994;
  assign n5126 = n5011 & n5125;
  assign n5127 = n5123 & n5124;
  assign n5128 = n5121 & n5122;
  assign n5129 = n5119 & n5120;
  assign n5130 = n399 & n1899;
  assign n5131 = n3003 & n3800;
  assign n5132 = n3994 & n4224;
  assign n5133 = n5007 & ~n5082;
  assign n5134 = n5087 & n5133;
  assign n5135 = n5131 & n5132;
  assign n5136 = n5129 & n5130;
  assign n5137 = n5127 & n5128;
  assign n5138 = n882 & n5126;
  assign n5139 = n2970 & n3627;
  assign n5140 = n5090 & n5139;
  assign n5141 = n5137 & n5138;
  assign n5142 = n5135 & n5136;
  assign n5143 = n4928 & n5134;
  assign n5144 = n4975 & n5040;
  assign n5145 = ~n5042 & n5144;
  assign n5146 = n5142 & n5143;
  assign n5147 = n5140 & n5141;
  assign n5148 = n5146 & n5147;
  assign n5149 = n5079 & n5145;
  assign n5150 = n5148 & n5149;
  assign po042 = ~n4380 | ~n5150;
  assign n5152 = ~n1153 & n4420;
  assign n5153 = n4388 & ~n5152;
  assign n5154 = n1898 & n5007;
  assign n5155 = n2095 & n5090;
  assign n5156 = ~n5153 & n5154;
  assign po043 = ~n5155 | ~n5156;
  assign n5158 = ~n4204 & n4207;
  assign n5159 = n2486 & n5158;
  assign n5160 = n329 & ~n5159;
  assign n5161 = n692 & n4059;
  assign n5162 = n2763 & n2781;
  assign n5163 = n4074 & n5056;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~pi027 & ~n5164;
  assign n5166 = pi013 & n3368;
  assign n5167 = ~n2594 & ~n5166;
  assign n5168 = ~n332 & ~n5167;
  assign n5169 = n4167 & ~n4189;
  assign n5170 = n5025 & n5169;
  assign n5171 = ~pi029 & n3031;
  assign n5172 = n1480 & n5171;
  assign n5173 = n902 & n4833;
  assign n5174 = n1326 & ~n4916;
  assign n5175 = ~n1033 & ~n1752;
  assign n5176 = ~n2597 & n5175;
  assign n5177 = ~n4820 & ~n5176;
  assign n5178 = n1753 & n5177;
  assign n5179 = n439 & n3473;
  assign n5180 = n1724 & ~n3060;
  assign n5181 = ~n2488 & n5180;
  assign n5182 = ~pi029 & n4830;
  assign n5183 = ~n1752 & n4125;
  assign n5184 = n3295 & ~n5183;
  assign n5185 = n960 & n1669;
  assign n5186 = n1325 & n5185;
  assign n5187 = n492 & n4203;
  assign n5188 = pi015 & n4047;
  assign n5189 = n2065 & n4970;
  assign n5190 = n1991 & ~n2522;
  assign n5191 = n1702 & ~n5190;
  assign n5192 = n4841 & ~n5191;
  assign n5193 = ~n4147 & n5192;
  assign n5194 = ~n1987 & ~n3167;
  assign n5195 = ~n5182 & n5194;
  assign n5196 = n4838 & n5195;
  assign n5197 = ~n5179 & ~n5181;
  assign n5198 = ~n5184 & ~n5186;
  assign n5199 = ~n5187 & n5198;
  assign n5200 = n5196 & n5197;
  assign n5201 = n2716 & ~n2909;
  assign n5202 = ~n3156 & n5029;
  assign n5203 = ~n5161 & ~n5172;
  assign n5204 = ~n5173 & ~n5178;
  assign n5205 = n5203 & n5204;
  assign n5206 = n5201 & n5202;
  assign n5207 = n5199 & n5200;
  assign n5208 = ~n5174 & n5207;
  assign n5209 = n5205 & n5206;
  assign n5210 = ~n3112 & n3796;
  assign n5211 = ~n3831 & ~n5165;
  assign n5212 = ~n5168 & n5170;
  assign n5213 = ~n5188 & n5212;
  assign n5214 = n5210 & n5211;
  assign n5215 = n5208 & n5209;
  assign n5216 = n4100 & n5215;
  assign n5217 = n5213 & n5214;
  assign n5218 = ~n4179 & n5217;
  assign n5219 = n4630 & n5216;
  assign n5220 = ~n5160 & n5189;
  assign n5221 = n5193 & n5220;
  assign n5222 = n5218 & n5219;
  assign po044 = ~n5221 | ~n5222;
  assign n5224 = ~n360 & n491;
  assign n5225 = ~n2779 & n5224;
  assign n5226 = n1336 & ~n1593;
  assign n5227 = n771 & n906;
  assign n5228 = n311 & n687;
  assign n5229 = ~n3075 & ~n5228;
  assign n5230 = n529 & ~n5229;
  assign n5231 = n2066 & n4138;
  assign n5232 = ~pi056 & n798;
  assign n5233 = n1513 & n5232;
  assign n5234 = pi061 & n5233;
  assign n5235 = ~n2707 & ~n2792;
  assign n5236 = n503 & ~n5235;
  assign n5237 = ~n790 & ~n1328;
  assign n5238 = pi029 & ~n5237;
  assign n5239 = ~n470 & ~n3872;
  assign n5240 = ~n5238 & n5239;
  assign n5241 = n329 & ~n5240;
  assign n5242 = n329 & ~n4495;
  assign n5243 = ~n1262 & ~n1482;
  assign n5244 = ~n1478 & n5243;
  assign n5245 = n5171 & ~n5244;
  assign n5246 = ~n2053 & n2744;
  assign n5247 = n1462 & ~n5246;
  assign n5248 = ~pi122 & n1279;
  assign n5249 = pi018 & n1277;
  assign n5250 = n345 & n5249;
  assign n5251 = ~pi122 & n1277;
  assign n5252 = n566 & n5251;
  assign n5253 = ~n5250 & ~n5252;
  assign n5254 = ~n5248 & n5253;
  assign n5255 = ~n3215 & ~n5012;
  assign n5256 = n5254 & n5255;
  assign n5257 = n750 & ~n1583;
  assign n5258 = n3103 & ~n5257;
  assign n5259 = n2746 & n4261;
  assign n5260 = n798 & n1583;
  assign n5261 = ~pi055 & pi056;
  assign n5262 = pi122 & n5261;
  assign n5263 = n2036 & n5262;
  assign n5264 = n3042 & n4213;
  assign n5265 = n2803 & n2929;
  assign n5266 = ~n2788 & n5265;
  assign n5267 = n5264 & n5266;
  assign n5268 = n791 & n2879;
  assign n5269 = n1891 & ~n5268;
  assign n5270 = n480 & n3979;
  assign n5271 = n3707 & ~n5270;
  assign n5272 = n492 & ~n5271;
  assign n5273 = n1338 & ~n2573;
  assign n5274 = n5040 & ~n5273;
  assign n5275 = ~n2590 & ~n5231;
  assign n5276 = ~n3115 & n5275;
  assign n5277 = ~n5230 & n5276;
  assign n5278 = ~n1133 & ~n3338;
  assign n5279 = ~n4238 & ~n5234;
  assign n5280 = ~n5247 & ~n5260;
  assign n5281 = ~n5263 & n5280;
  assign n5282 = n5278 & n5279;
  assign n5283 = ~n3976 & n5277;
  assign n5284 = ~n4752 & ~n4852;
  assign n5285 = ~n5236 & ~n5258;
  assign n5286 = n5284 & n5285;
  assign n5287 = n5282 & n5283;
  assign n5288 = n342 & n5281;
  assign n5289 = n595 & ~n5259;
  assign n5290 = n5288 & n5289;
  assign n5291 = n5286 & n5287;
  assign n5292 = n871 & n2762;
  assign n5293 = ~n3049 & ~n3527;
  assign n5294 = n3986 & n4921;
  assign n5295 = n5293 & n5294;
  assign n5296 = n5291 & n5292;
  assign n5297 = n1043 & n5290;
  assign n5298 = n3729 & ~n4219;
  assign n5299 = ~n5225 & ~n5226;
  assign n5300 = ~n5241 & n5299;
  assign n5301 = n5297 & n5298;
  assign n5302 = n5295 & n5296;
  assign n5303 = n806 & n4185;
  assign n5304 = ~n5227 & ~n5242;
  assign n5305 = ~n5245 & n5256;
  assign n5306 = n5304 & n5305;
  assign n5307 = n5302 & n5303;
  assign n5308 = n5300 & n5301;
  assign n5309 = n881 & ~n2468;
  assign n5310 = n2617 & n3174;
  assign n5311 = n3626 & n4115;
  assign n5312 = n5269 & ~n5272;
  assign n5313 = n5311 & n5312;
  assign n5314 = n5309 & n5310;
  assign n5315 = n5307 & n5308;
  assign n5316 = n5306 & n5315;
  assign n5317 = n5313 & n5314;
  assign n5318 = n5316 & n5317;
  assign n5319 = n5267 & n5274;
  assign n5320 = n5318 & n5319;
  assign n5321 = n3006 & n5079;
  assign n5322 = n5320 & n5321;
  assign po046 = ~n4382 | ~n5322;
  assign n5324 = ~n2902 & ~n3542;
  assign n5325 = ~n1328 & ~n1335;
  assign n5326 = n740 & ~n5325;
  assign n5327 = ~n1518 & n2745;
  assign n5328 = pi027 & n2763;
  assign n5329 = ~n2782 & n5328;
  assign n5330 = ~n360 & n1241;
  assign n5331 = n3068 & n5330;
  assign n5332 = ~n2724 & ~n3832;
  assign n5333 = n329 & ~n5332;
  assign n5334 = ~n3365 & ~n5333;
  assign n5335 = ~n3033 & n5334;
  assign n5336 = pi029 & ~n5335;
  assign n5337 = ~n990 & n3814;
  assign n5338 = ~n2409 & ~n3545;
  assign n5339 = ~n5327 & n5338;
  assign n5340 = ~n2661 & ~n2670;
  assign n5341 = ~n4175 & n5324;
  assign n5342 = ~n5331 & n5341;
  assign n5343 = n5339 & n5340;
  assign n5344 = ~n5000 & ~n5337;
  assign n5345 = n5343 & n5344;
  assign n5346 = ~n4101 & n5342;
  assign n5347 = n4920 & ~n5326;
  assign n5348 = n5346 & n5347;
  assign n5349 = n4981 & n5345;
  assign n5350 = ~n5329 & n5349;
  assign n5351 = ~n3292 & n5348;
  assign n5352 = n5350 & n5351;
  assign n5353 = n3725 & n5352;
  assign po047 = n5336 | ~n5353;
  assign n5355 = ~n864 & ~n1572;
  assign po050 = ~n3792 | ~n5355;
  assign n5357 = ~n3887 & ~n4073;
  assign n5358 = n308 & n349;
  assign n5359 = ~pi028 & pi039;
  assign n5360 = n311 & ~n5359;
  assign n5361 = n802 & n5360;
  assign n5362 = n5358 & n5361;
  assign n5363 = n307 & n492;
  assign n5364 = n759 & n5363;
  assign n5365 = ~n5362 & ~n5364;
  assign n5366 = pi108 & ~n5365;
  assign n5367 = n1539 & n2835;
  assign n5368 = n2381 & n5367;
  assign n5369 = ~n466 & ~n622;
  assign n5370 = n2597 & ~n5369;
  assign n5371 = n460 & n1776;
  assign n5372 = n573 & n598;
  assign n5373 = n569 & n5372;
  assign n5374 = ~pi029 & n3818;
  assign n5375 = n580 & n1795;
  assign n5376 = n466 & n5375;
  assign n5377 = pi009 & n3898;
  assign n5378 = ~pi039 & n992;
  assign n5379 = n405 & n1922;
  assign n5380 = n5378 & n5379;
  assign n5381 = n417 & n1049;
  assign n5382 = ~n2938 & ~n5381;
  assign n5383 = n293 & n1355;
  assign n5384 = ~n5382 & n5383;
  assign n5385 = n329 & ~n780;
  assign n5386 = n499 & n4827;
  assign n5387 = n606 & n1697;
  assign n5388 = ~n1675 & ~n5387;
  assign n5389 = n960 & ~n5388;
  assign n5390 = ~pi108 & n760;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = n492 & ~n5391;
  assign n5393 = ~pi039 & n492;
  assign n5394 = n751 & n1053;
  assign n5395 = n5393 & n5394;
  assign n5396 = n2487 & n3331;
  assign n5397 = n315 & n758;
  assign n5398 = ~n3203 & n5397;
  assign n5399 = ~pi019 & n2484;
  assign n5400 = ~n3855 & ~n5399;
  assign n5401 = n626 & ~n1752;
  assign n5402 = n628 & ~n5401;
  assign n5403 = n995 & n5393;
  assign n5404 = ~n5402 & ~n5403;
  assign n5405 = n798 & n1435;
  assign n5406 = ~n2660 & ~n5405;
  assign n5407 = n449 & ~n1006;
  assign n5408 = n371 & n5407;
  assign n5409 = ~n2651 & ~n5408;
  assign n5410 = n5406 & n5409;
  assign n5411 = n4385 & ~n5410;
  assign n5412 = ~pi045 & n336;
  assign n5413 = n1523 & n5412;
  assign n5414 = n599 & n5413;
  assign n5415 = ~n5411 & ~n5414;
  assign n5416 = ~pi045 & n2844;
  assign n5417 = ~n1228 & ~n2692;
  assign n5418 = n1092 & ~n5417;
  assign n5419 = n330 & n2791;
  assign n5420 = n2410 & ~n5419;
  assign n5421 = ~n5418 & n5420;
  assign n5422 = n5087 & n5421;
  assign n5423 = n646 & ~n3039;
  assign n5424 = ~pi122 & ~n4625;
  assign n5425 = ~n381 & n383;
  assign n5426 = ~n2873 & ~n3594;
  assign n5427 = ~n2093 & n5426;
  assign n5428 = ~n3740 & n5427;
  assign n5429 = n2311 & n5428;
  assign n5430 = ~n5423 & ~n5424;
  assign n5431 = n5429 & n5430;
  assign n5432 = ~n5425 & n5431;
  assign n5433 = ~pi039 & ~n5432;
  assign n5434 = ~n1790 & ~n2623;
  assign n5435 = n303 & ~n5434;
  assign n5436 = ~n1481 & n3031;
  assign n5437 = n294 & n532;
  assign n5438 = ~n350 & ~n452;
  assign n5439 = ~pi004 & ~n5438;
  assign n5440 = ~n479 & n747;
  assign n5441 = ~pi001 & ~pi006;
  assign n5442 = ~pi003 & ~n5441;
  assign n5443 = ~n5440 & n5442;
  assign n5444 = ~n5439 & ~n5443;
  assign n5445 = ~pi017 & ~n3639;
  assign n5446 = ~pi018 & ~n5445;
  assign n5447 = pi016 & ~n5446;
  assign n5448 = n350 & ~n5447;
  assign n5449 = n292 & n5448;
  assign n5450 = n5444 & ~n5449;
  assign n5451 = ~pi056 & ~n5450;
  assign n5452 = n293 & n4029;
  assign n5453 = ~n321 & n606;
  assign n5454 = ~n702 & ~n5453;
  assign n5455 = pi008 & n607;
  assign n5456 = ~n5454 & n5455;
  assign n5457 = ~pi008 & pi009;
  assign n5458 = ~n1782 & n5457;
  assign n5459 = ~n5456 & ~n5458;
  assign n5460 = n5452 & ~n5459;
  assign n5461 = ~pi003 & n5441;
  assign n5462 = n1708 & n2695;
  assign n5463 = n416 & n5462;
  assign n5464 = n350 & n5463;
  assign n5465 = ~n455 & ~n5461;
  assign n5466 = ~n5464 & n5465;
  assign n5467 = ~n5460 & n5466;
  assign n5468 = ~n5451 & n5467;
  assign n5469 = n5437 & ~n5468;
  assign n5470 = ~pi000 & n532;
  assign n5471 = pi002 & ~n970;
  assign n5472 = pi000 & ~n5471;
  assign n5473 = ~pi056 & n5472;
  assign n5474 = n532 & n5473;
  assign n5475 = ~n5470 & ~n5474;
  assign n5476 = ~n5469 & n5475;
  assign n5477 = n1228 & ~n5476;
  assign n5478 = ~n5436 & ~n5477;
  assign n5479 = n1660 & n1742;
  assign n5480 = ~n1501 & ~n2357;
  assign n5481 = ~n2578 & ~n5479;
  assign n5482 = n5480 & n5481;
  assign n5483 = n492 & ~n5482;
  assign n5484 = n780 & ~n797;
  assign n5485 = n798 & ~n5484;
  assign n5486 = n587 & n2716;
  assign n5487 = n740 & ~n991;
  assign n5488 = ~n828 & n5487;
  assign n5489 = ~pi045 & ~n1354;
  assign n5490 = ~pi039 & n5489;
  assign n5491 = n812 & ~n3009;
  assign n5492 = n347 & n5491;
  assign n5493 = n405 & n827;
  assign n5494 = ~pi122 & ~n3009;
  assign n5495 = n5493 & n5494;
  assign n5496 = ~n1309 & ~n2880;
  assign n5497 = n1465 & n5496;
  assign n5498 = ~n5495 & n5497;
  assign n5499 = ~pi045 & ~n5498;
  assign n5500 = ~n5492 & ~n5499;
  assign n5501 = n330 & ~n5500;
  assign n5502 = ~n818 & ~n5493;
  assign n5503 = n330 & n4385;
  assign n5504 = ~n5502 & n5503;
  assign n5505 = ~pi023 & n1426;
  assign n5506 = ~n348 & ~n510;
  assign n5507 = n2229 & ~n5506;
  assign n5508 = n949 & n2251;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~n5505 & n5509;
  assign n5511 = n2381 & ~n5510;
  assign n5512 = ~n5504 & ~n5511;
  assign n5513 = ~n5490 & n5512;
  assign n5514 = ~n5501 & n5513;
  assign n5515 = ~n2232 & n2233;
  assign n5516 = n1507 & ~n2979;
  assign n5517 = ~n5515 & n5516;
  assign n5518 = ~n2246 & n5517;
  assign n5519 = n453 & n2932;
  assign n5520 = ~n2974 & ~n5519;
  assign n5521 = ~n1420 & ~n3046;
  assign n5522 = ~n1394 & n5521;
  assign n5523 = n5520 & n5522;
  assign n5524 = ~n2302 & ~n2330;
  assign n5525 = n5523 & n5524;
  assign n5526 = n5518 & n5525;
  assign n5527 = ~n474 & ~n5526;
  assign n5528 = n417 & n599;
  assign n5529 = n1078 & ~n5528;
  assign n5530 = n293 & ~n5529;
  assign n5531 = ~n2243 & n2995;
  assign n5532 = ~n5530 & n5531;
  assign n5533 = n345 & ~n5532;
  assign n5534 = ~n873 & ~n5533;
  assign n5535 = ~n5527 & n5534;
  assign n5536 = ~pi039 & ~n5535;
  assign n5537 = n752 & ~n828;
  assign n5538 = ~n740 & ~n5393;
  assign n5539 = n5537 & ~n5538;
  assign n5540 = pi045 & ~n831;
  assign n5541 = ~n828 & ~n5540;
  assign n5542 = n879 & ~n5541;
  assign n5543 = n492 & ~n820;
  assign n5544 = ~pi044 & n473;
  assign n5545 = pi122 & ~n5544;
  assign n5546 = ~pi005 & ~n5545;
  assign n5547 = pi022 & n3621;
  assign n5548 = ~n1388 & ~n2256;
  assign n5549 = ~n5547 & n5548;
  assign n5550 = n336 & n5546;
  assign n5551 = ~n5549 & n5550;
  assign n5552 = ~n934 & ~n1060;
  assign n5553 = ~n2255 & n5552;
  assign n5554 = n510 & n930;
  assign n5555 = ~n3071 & n5553;
  assign n5556 = ~n5554 & n5555;
  assign n5557 = n3092 & n5556;
  assign n5558 = ~pi022 & n1722;
  assign n5559 = n412 & n492;
  assign n5560 = pi022 & ~n2951;
  assign n5561 = ~n1259 & ~n5558;
  assign n5562 = ~n5559 & n5561;
  assign n5563 = ~n5560 & n5562;
  assign n5564 = ~n2258 & n5563;
  assign n5565 = n5557 & n5564;
  assign n5566 = n361 & ~n5565;
  assign n5567 = ~n5542 & ~n5551;
  assign n5568 = ~n5543 & n5567;
  assign n5569 = ~n5566 & n5568;
  assign n5570 = ~pi039 & ~n5569;
  assign n5571 = n791 & ~n2773;
  assign n5572 = ~n2669 & ~n3637;
  assign n5573 = ~n807 & ~n2539;
  assign n5574 = n5572 & n5573;
  assign n5575 = n1376 & ~n5574;
  assign n5576 = n353 & n568;
  assign n5577 = ~n5547 & ~n5576;
  assign n5578 = n293 & ~n5577;
  assign n5579 = n518 & n971;
  assign n5580 = n306 & n2264;
  assign n5581 = ~n2291 & ~n5579;
  assign n5582 = ~n5580 & n5581;
  assign n5583 = ~n5578 & n5582;
  assign n5584 = n4385 & ~n5583;
  assign n5585 = n1397 & n4826;
  assign n5586 = ~n5571 & ~n5585;
  assign n5587 = ~n5575 & n5586;
  assign n5588 = ~n5584 & n5587;
  assign n5589 = ~pi039 & ~n5588;
  assign n5590 = ~n1897 & ~n2105;
  assign n5591 = ~n1169 & n5590;
  assign n5592 = ~pi056 & ~n5591;
  assign n5593 = ~pi056 & ~pi122;
  assign n5594 = pi044 & ~pi055;
  assign n5595 = pi045 & n5594;
  assign n5596 = n1134 & ~n5595;
  assign n5597 = ~n5593 & ~n5596;
  assign n5598 = n2858 & ~n4417;
  assign n5599 = n5596 & ~n5598;
  assign n5600 = n2864 & ~n5599;
  assign n5601 = ~n5597 & ~n5600;
  assign n5602 = n4391 & n4410;
  assign n5603 = ~pi056 & ~n5602;
  assign n5604 = ~pi045 & n306;
  assign n5605 = n4398 & n5604;
  assign n5606 = n1215 & n5593;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = ~n5603 & n5607;
  assign n5609 = ~n5592 & n5608;
  assign n5610 = ~n5601 & n5609;
  assign n5611 = n1517 & n3637;
  assign n5612 = n603 & n866;
  assign n5613 = ~n5363 & ~n5546;
  assign n5614 = ~pi004 & ~n5613;
  assign n5615 = ~n1357 & ~n1620;
  assign n5616 = ~n360 & ~n5615;
  assign n5617 = ~n5614 & ~n5616;
  assign n5618 = n3979 & ~n5617;
  assign n5619 = ~n3011 & ~n4385;
  assign n5620 = pi001 & ~pi005;
  assign n5621 = n4385 & ~n5620;
  assign n5622 = n311 & ~n5621;
  assign n5623 = ~n5619 & n5622;
  assign n5624 = n751 & ~n5545;
  assign n5625 = pi004 & n4385;
  assign n5626 = n2932 & n5625;
  assign n5627 = ~n5624 & ~n5626;
  assign n5628 = n292 & ~n5627;
  assign n5629 = n349 & n5544;
  assign n5630 = n5379 & n5629;
  assign n5631 = ~pi029 & n3012;
  assign n5632 = ~n633 & ~n2297;
  assign n5633 = n1922 & n2932;
  assign n5634 = n5632 & ~n5633;
  assign n5635 = ~n5545 & ~n5634;
  assign n5636 = n2341 & ~n5630;
  assign n5637 = ~n5623 & ~n5631;
  assign n5638 = n5636 & n5637;
  assign n5639 = ~n5628 & ~n5635;
  assign n5640 = n5638 & n5639;
  assign n5641 = ~pi039 & ~n5640;
  assign n5642 = n1355 & n2774;
  assign n5643 = ~n755 & ~n1623;
  assign n5644 = ~n5642 & n5643;
  assign n5645 = n492 & ~n5644;
  assign n5646 = ~n5611 & ~n5612;
  assign n5647 = ~n5618 & ~n5645;
  assign n5648 = n5646 & n5647;
  assign n5649 = ~n5641 & n5648;
  assign n5650 = n851 & n5649;
  assign n5651 = n4433 & n5650;
  assign n5652 = ~n5589 & n5651;
  assign n5653 = n5610 & n5652;
  assign n5654 = ~n5570 & n5653;
  assign n5655 = ~n5539 & n5654;
  assign n5656 = ~n2396 & ~n2916;
  assign n5657 = ~n2883 & n5656;
  assign n5658 = n2238 & n5657;
  assign n5659 = n3065 & n5658;
  assign n5660 = ~pi045 & ~n5659;
  assign n5661 = ~pi056 & n1530;
  assign n5662 = n1249 & ~n5661;
  assign n5663 = n3025 & n5662;
  assign n5664 = n2646 & ~n5663;
  assign n5665 = n330 & n1468;
  assign n5666 = ~n1444 & ~n2395;
  assign n5667 = ~n2992 & n5666;
  assign n5668 = ~n990 & n1461;
  assign n5669 = n293 & n5668;
  assign n5670 = n5667 & ~n5669;
  assign n5671 = ~n5665 & n5670;
  assign n5672 = ~n2718 & n5671;
  assign n5673 = ~n2805 & n5672;
  assign n5674 = ~pi045 & ~n5673;
  assign n5675 = n2648 & ~n5674;
  assign n5676 = ~n1177 & n2828;
  assign n5677 = n572 & n2365;
  assign n5678 = ~n5676 & n5677;
  assign n5679 = n1029 & n1228;
  assign n5680 = n330 & n1440;
  assign n5681 = ~n2393 & ~n5680;
  assign n5682 = ~n5679 & n5681;
  assign n5683 = n2272 & ~n2281;
  assign n5684 = n416 & ~n5683;
  assign n5685 = ~n1028 & n3020;
  assign n5686 = n572 & ~n5685;
  assign n5687 = n5682 & ~n5686;
  assign n5688 = ~n5684 & n5687;
  assign n5689 = ~pi045 & ~n5688;
  assign n5690 = n453 & n1177;
  assign n5691 = ~n1920 & n2894;
  assign n5692 = n2686 & ~n5690;
  assign n5693 = n4544 & n5692;
  assign n5694 = n5691 & n5693;
  assign n5695 = n4427 & ~n5694;
  assign n5696 = ~n5664 & ~n5678;
  assign n5697 = n5675 & n5696;
  assign n5698 = ~n5689 & n5697;
  assign n5699 = ~n5660 & n5698;
  assign n5700 = ~n5695 & n5699;
  assign n5701 = n492 & n1435;
  assign n5702 = n1134 & n5701;
  assign n5703 = n330 & ~n2900;
  assign n5704 = ~n2755 & ~n3768;
  assign n5705 = ~n5703 & n5704;
  assign n5706 = ~pi056 & ~n5705;
  assign n5707 = ~pi056 & n492;
  assign n5708 = ~n3113 & n5707;
  assign n5709 = ~n5702 & ~n5708;
  assign n5710 = ~n5706 & n5709;
  assign n5711 = n5700 & n5710;
  assign n5712 = n2381 & n2848;
  assign n5713 = n5711 & ~n5712;
  assign n5714 = ~n2060 & ~n5380;
  assign n5715 = ~n4961 & ~n5386;
  assign n5716 = ~n5395 & n5715;
  assign n5717 = ~n432 & n5714;
  assign n5718 = ~n3183 & ~n5373;
  assign n5719 = ~n5376 & ~n5377;
  assign n5720 = ~n5396 & ~n5398;
  assign n5721 = n5719 & n5720;
  assign n5722 = n5717 & n5718;
  assign n5723 = ~n2370 & n5716;
  assign n5724 = ~n3270 & ~n4164;
  assign n5725 = ~n4415 & n5357;
  assign n5726 = n5724 & n5725;
  assign n5727 = n5722 & n5723;
  assign n5728 = ~n5366 & n5721;
  assign n5729 = ~n5368 & ~n5370;
  assign n5730 = ~n5371 & ~n5374;
  assign n5731 = n5400 & n5404;
  assign n5732 = n5730 & n5731;
  assign n5733 = n5728 & n5729;
  assign n5734 = n5726 & n5727;
  assign n5735 = ~n5384 & ~n5385;
  assign n5736 = ~n5392 & n5486;
  assign n5737 = ~n5488 & n5736;
  assign n5738 = n5734 & n5735;
  assign n5739 = n5732 & n5733;
  assign n5740 = ~n5435 & ~n5483;
  assign n5741 = ~n5485 & n5740;
  assign n5742 = n5738 & n5739;
  assign n5743 = n3298 & n5737;
  assign n5744 = n3914 & n5415;
  assign n5745 = ~n5416 & n5744;
  assign n5746 = n5742 & n5743;
  assign n5747 = n5478 & n5741;
  assign n5748 = n5746 & n5747;
  assign n5749 = n4384 & n5745;
  assign n5750 = n5422 & ~n5433;
  assign n5751 = n5749 & n5750;
  assign n5752 = n5514 & n5748;
  assign n5753 = n5751 & n5752;
  assign n5754 = ~n5536 & n5753;
  assign n5755 = n5655 & n5754;
  assign po052 = ~n5713 | ~n5755;
  assign n5757 = n2365 & ~n2779;
  assign n5758 = ~n1755 & ~n5757;
  assign n5759 = ~n2594 & n5193;
  assign n5760 = ~n3163 & ~n4048;
  assign n5761 = n329 & ~n783;
  assign n5762 = ~n5085 & ~n5761;
  assign n5763 = n1620 & n2792;
  assign n5764 = ~n3294 & ~n5763;
  assign n5765 = ~n408 & ~n2692;
  assign n5766 = n1092 & ~n5765;
  assign n5767 = ~n622 & ~n4059;
  assign n5768 = n1702 & ~n5767;
  assign n5769 = ~n2943 & n5267;
  assign n5770 = ~pi039 & ~n5769;
  assign n5771 = n5517 & n5523;
  assign n5772 = n1355 & ~n5771;
  assign n5773 = ~pi039 & n873;
  assign n5774 = pi034 & n5397;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = ~pi039 & n345;
  assign n5777 = ~n378 & ~n2330;
  assign n5778 = n2990 & n5777;
  assign n5779 = n2997 & n5778;
  assign n5780 = n5776 & ~n5779;
  assign n5781 = n2511 & ~n3620;
  assign n5782 = n573 & ~n2827;
  assign n5783 = ~n2326 & ~n5379;
  assign n5784 = n5378 & ~n5783;
  assign n5785 = n349 & ~n3224;
  assign n5786 = n1586 & n5785;
  assign n5787 = ~n1585 & n5786;
  assign n5788 = ~n429 & ~n4492;
  assign n5789 = n1523 & ~n5788;
  assign n5790 = ~n799 & n2774;
  assign n5791 = ~n5784 & ~n5790;
  assign n5792 = ~n5364 & n5791;
  assign n5793 = ~n5787 & n5792;
  assign n5794 = n2377 & n5793;
  assign n5795 = ~n5789 & n5794;
  assign n5796 = n588 & n2372;
  assign n5797 = ~n5782 & n5796;
  assign n5798 = ~n5781 & n5795;
  assign n5799 = n5797 & n5798;
  assign n5800 = n5775 & n5799;
  assign n5801 = ~n5780 & n5800;
  assign n5802 = ~n5772 & n5801;
  assign n5803 = ~n5770 & n5802;
  assign n5804 = pi029 & n1502;
  assign n5805 = ~n3237 & ~n3527;
  assign n5806 = ~n5804 & n5805;
  assign n5807 = ~n1841 & n5806;
  assign n5808 = ~n4811 & n5807;
  assign n5809 = n4206 & n4931;
  assign n5810 = n471 & n5809;
  assign n5811 = n492 & ~n5810;
  assign n5812 = pi002 & n5461;
  assign n5813 = pi000 & ~n5812;
  assign n5814 = ~n534 & ~n5813;
  assign n5815 = pi000 & ~n534;
  assign n5816 = pi002 & n5815;
  assign n5817 = n350 & n5816;
  assign n5818 = n5463 & n5817;
  assign n5819 = ~n5814 & ~n5818;
  assign n5820 = ~n2614 & ~n5819;
  assign n5821 = n416 & n5448;
  assign n5822 = n5444 & ~n5821;
  assign n5823 = ~pi056 & ~n5822;
  assign n5824 = ~n455 & ~n5460;
  assign n5825 = ~n5823 & n5824;
  assign n5826 = n294 & ~n5825;
  assign n5827 = ~n5473 & ~n5826;
  assign n5828 = ~n534 & n798;
  assign n5829 = ~n5827 & n5828;
  assign n5830 = n293 & n5817;
  assign n5831 = n452 & n5816;
  assign n5832 = n549 & n5831;
  assign n5833 = ~n5830 & ~n5832;
  assign n5834 = n5393 & ~n5833;
  assign n5835 = ~pi002 & n5815;
  assign n5836 = pi001 & n1338;
  assign n5837 = n970 & ~n1400;
  assign n5838 = ~pi006 & n318;
  assign n5839 = n322 & n5838;
  assign n5840 = ~n5837 & ~n5839;
  assign n5841 = n518 & n740;
  assign n5842 = ~n5840 & n5841;
  assign n5843 = ~n5836 & ~n5842;
  assign n5844 = n5835 & ~n5843;
  assign n5845 = ~n5820 & ~n5834;
  assign n5846 = ~n5844 & n5845;
  assign n5847 = ~n5829 & n5846;
  assign n5848 = n3331 & n4094;
  assign n5849 = ~n722 & n2050;
  assign n5850 = ~n1784 & ~n5849;
  assign n5851 = n1787 & ~n5850;
  assign n5852 = ~n1718 & n2182;
  assign n5853 = n3295 & ~n5852;
  assign n5854 = ~n290 & ~n1670;
  assign n5855 = n1752 & ~n5854;
  assign n5856 = n960 & n5855;
  assign n5857 = n492 & n1746;
  assign n5858 = n2487 & n5857;
  assign n5859 = ~n3330 & ~n4912;
  assign n5860 = n1990 & ~n5859;
  assign n5861 = n290 & n438;
  assign n5862 = ~n5021 & n5861;
  assign n5863 = ~n5848 & ~n5856;
  assign n5864 = ~n5858 & n5863;
  assign n5865 = ~n5186 & ~n5853;
  assign n5866 = ~n5860 & ~n5862;
  assign n5867 = n5865 & n5866;
  assign n5868 = n4989 & n5864;
  assign n5869 = ~n5851 & n5868;
  assign n5870 = ~n4915 & n5867;
  assign n5871 = n5869 & n5870;
  assign n5872 = ~n1033 & ~n5056;
  assign n5873 = n2623 & ~n5872;
  assign n5874 = n1024 & n1674;
  assign n5875 = ~n994 & ~n5358;
  assign n5876 = n5361 & ~n5875;
  assign n5877 = n1264 & ~n5244;
  assign n5878 = n354 & n2512;
  assign n5879 = n482 & n3591;
  assign n5880 = ~n566 & n5879;
  assign n5881 = n421 & n3605;
  assign n5882 = ~n2513 & ~n2798;
  assign n5883 = n598 & ~n5882;
  assign n5884 = n596 & n1684;
  assign n5885 = n510 & n3580;
  assign n5886 = ~n3600 & ~n5885;
  assign n5887 = pi020 & n776;
  assign n5888 = ~n5886 & n5887;
  assign n5889 = ~n5883 & ~n5884;
  assign n5890 = ~n5888 & n5889;
  assign n5891 = n418 & ~n5890;
  assign n5892 = ~n410 & ~n668;
  assign n5893 = n3251 & ~n5892;
  assign n5894 = ~n4621 & ~n5878;
  assign n5895 = ~n5880 & ~n5881;
  assign n5896 = n5894 & n5895;
  assign n5897 = ~n5891 & ~n5893;
  assign n5898 = n5896 & n5897;
  assign n5899 = pi029 & n2781;
  assign n5900 = pi027 & n5899;
  assign n5901 = ~n5273 & ~n5900;
  assign n5902 = ~n2621 & n5898;
  assign n5903 = ~n5877 & n5902;
  assign n5904 = n4857 & n5903;
  assign n5905 = n5901 & n5904;
  assign n5906 = n4928 & n5905;
  assign n5907 = ~n1588 & ~n3234;
  assign n5908 = ~n5876 & n5907;
  assign n5909 = ~n3183 & n5908;
  assign n5910 = ~n1045 & n5909;
  assign n5911 = n686 & n4775;
  assign n5912 = ~n5487 & ~n5874;
  assign n5913 = n5911 & n5912;
  assign n5914 = n2070 & n5910;
  assign n5915 = n5764 & ~n5766;
  assign n5916 = ~n5768 & ~n5873;
  assign n5917 = n5915 & n5916;
  assign n5918 = n5913 & n5914;
  assign n5919 = n1622 & ~n5010;
  assign n5920 = n5420 & n5919;
  assign n5921 = n5917 & n5918;
  assign n5922 = n1251 & n4078;
  assign n5923 = n4602 & n4967;
  assign n5924 = n5083 & n5256;
  assign n5925 = n5758 & n5760;
  assign n5926 = n5762 & n5871;
  assign n5927 = n5925 & n5926;
  assign n5928 = n5923 & n5924;
  assign n5929 = n5921 & n5922;
  assign n5930 = ~n5811 & n5920;
  assign n5931 = n5847 & n5930;
  assign n5932 = n5928 & n5929;
  assign n5933 = n5808 & n5927;
  assign n5934 = n5932 & n5933;
  assign n5935 = n5040 & n5931;
  assign n5936 = n5759 & n5935;
  assign n5937 = n5906 & n5934;
  assign n5938 = n5936 & n5937;
  assign n5939 = n5655 & n5938;
  assign po053 = ~n5803 | ~n5939;
  assign n5941 = pi002 & n1355;
  assign n5942 = n378 & n5941;
  assign n5943 = pi019 & po025;
  assign n5944 = ~n2996 & ~n4037;
  assign n5945 = n5776 & ~n5944;
  assign n5946 = n938 & n5367;
  assign n5947 = ~n2851 & ~n5946;
  assign n5948 = n5514 & n5947;
  assign n5949 = n5415 & n5948;
  assign po157 = ~n5711 | ~n5949;
  assign n5951 = ~n555 & ~n5757;
  assign n5952 = ~n393 & ~n2042;
  assign n5953 = ~n557 & ~n2332;
  assign n5954 = ~n3543 & n5953;
  assign n5955 = n5952 & n5954;
  assign n5956 = n4273 & n5955;
  assign n5957 = ~pi039 & ~n5956;
  assign n5958 = ~n3999 & ~n5942;
  assign n5959 = ~n5786 & n5958;
  assign n5960 = n2591 & n5959;
  assign n5961 = ~n5804 & n5960;
  assign n5962 = ~n5943 & ~n5945;
  assign n5963 = n5961 & n5962;
  assign n5964 = n5951 & n5963;
  assign n5965 = ~n5957 & n5964;
  assign n5966 = n5847 & n5965;
  assign po054 = po157 | ~n5966;
  assign n5968 = n1011 & n5861;
  assign n5969 = ~n781 & ~n2774;
  assign n5970 = n798 & ~n5969;
  assign n5971 = ~n782 & ~n3277;
  assign n5972 = ~n1583 & n5971;
  assign n5973 = n330 & ~n5972;
  assign n5974 = n780 & ~n5970;
  assign n5975 = ~n5973 & n5974;
  assign n5976 = ~n799 & ~n5975;
  assign n5977 = n740 & ~n4044;
  assign n5978 = n5764 & ~n5977;
  assign n5979 = ~n5976 & n5978;
  assign n5980 = n5422 & n5979;
  assign n5981 = n2486 & n4205;
  assign n5982 = n492 & ~n5981;
  assign n5983 = ~n5858 & ~n5873;
  assign n5984 = ~pi011 & ~n5983;
  assign n5985 = ~n510 & n3269;
  assign n5986 = n4051 & ~n5985;
  assign n5987 = ~pi023 & n3617;
  assign n5988 = n3619 & ~n5987;
  assign n5989 = n2511 & ~n5988;
  assign n5990 = ~n4123 & n5185;
  assign n5991 = ~n2371 & ~n5990;
  assign n5992 = n4802 & n5991;
  assign n5993 = n1989 & n1990;
  assign n5994 = pi016 & n2512;
  assign n5995 = ~n3053 & ~n5994;
  assign n5996 = n486 & ~n5995;
  assign n5997 = ~n1705 & ~n4079;
  assign n5998 = ~pi013 & ~n5997;
  assign n5999 = n368 & n3295;
  assign n6000 = ~n5008 & ~n5996;
  assign n6001 = ~n5968 & n6000;
  assign n6002 = ~n5993 & ~n5999;
  assign n6003 = n6001 & n6002;
  assign n6004 = ~n2575 & ~n3488;
  assign n6005 = ~n3590 & n4837;
  assign n6006 = ~n5998 & n6005;
  assign n6007 = n6003 & n6004;
  assign n6008 = ~n1755 & ~n2368;
  assign n6009 = n3572 & n6008;
  assign n6010 = n6006 & n6007;
  assign n6011 = ~n1250 & ~n1792;
  assign n6012 = n5986 & ~n5989;
  assign n6013 = n6011 & n6012;
  assign n6014 = n6009 & n6010;
  assign n6015 = ~n5984 & n6014;
  assign n6016 = n5192 & n6013;
  assign n6017 = n5807 & n6016;
  assign n6018 = ~n5982 & n6015;
  assign n6019 = n5992 & n6018;
  assign n6020 = n5980 & n6017;
  assign n6021 = n6019 & n6020;
  assign po055 = ~n5906 | ~n6021;
  assign n6023 = n2779 & ~n4067;
  assign n6024 = pi029 & ~n6023;
  assign n6025 = n2716 & n3546;
  assign n6026 = n5009 & n6025;
  assign n6027 = ~n5877 & n6026;
  assign n6028 = n5478 & n6027;
  assign n6029 = n5901 & ~n6024;
  assign n6030 = n6028 & n6029;
  assign n6031 = n5808 & n6030;
  assign n6032 = n5980 & n6031;
  assign po056 = po157 | ~n6032;
  assign n6034 = n1478 & n3031;
  assign n6035 = ~n1278 & ~n3054;
  assign n6036 = n2653 & n5406;
  assign n6037 = pi122 & ~n6036;
  assign n6038 = n6035 & ~n6037;
  assign n6039 = ~pi045 & ~n6038;
  assign n6040 = n492 & ~n4932;
  assign n6041 = pi060 & ~n1248;
  assign n6042 = n1250 & ~n6041;
  assign n6043 = n1790 & n4058;
  assign n6044 = n667 & n1531;
  assign n6045 = n5251 & n6044;
  assign n6046 = n372 & n1033;
  assign n6047 = ~n5249 & ~n6046;
  assign n6048 = n5544 & ~n6047;
  assign n6049 = n302 & n4385;
  assign n6050 = n372 & n6049;
  assign n6051 = ~n997 & ~n3172;
  assign n6052 = n5393 & ~n6051;
  assign n6053 = pi045 & n5252;
  assign n6054 = ~n368 & ~n606;
  assign n6055 = ~n1325 & ~n2029;
  assign n6056 = n6054 & n6055;
  assign n6057 = n439 & ~n6056;
  assign n6058 = ~n5027 & ~n6050;
  assign n6059 = ~n305 & n6058;
  assign n6060 = n1589 & ~n2054;
  assign n6061 = ~n4923 & ~n6052;
  assign n6062 = ~n6057 & n6061;
  assign n6063 = n6059 & n6060;
  assign n6064 = n3546 & n4072;
  assign n6065 = ~n4407 & n4775;
  assign n6066 = n5404 & ~n6045;
  assign n6067 = n6065 & n6066;
  assign n6068 = n6063 & n6064;
  assign n6069 = ~n1321 & n6062;
  assign n6070 = ~n4811 & ~n6034;
  assign n6071 = ~n6043 & ~n6048;
  assign n6072 = ~n6053 & n6071;
  assign n6073 = n6069 & n6070;
  assign n6074 = n6067 & n6068;
  assign n6075 = n5898 & n6074;
  assign n6076 = n6072 & n6073;
  assign n6077 = n5806 & n5951;
  assign n6078 = ~n6042 & n6077;
  assign n6079 = n6075 & n6076;
  assign n6080 = n3299 & ~n6039;
  assign n6081 = ~n6040 & n6080;
  assign n6082 = n6078 & n6079;
  assign n6083 = n6081 & n6082;
  assign n6084 = n4975 & n6083;
  assign n6085 = n5274 & n5948;
  assign n6086 = n6084 & n6085;
  assign n6087 = n5654 & n6086;
  assign n6088 = n5711 & n6087;
  assign po057 = ~n5803 | ~n6088;
  assign n6090 = ~n468 & n5809;
  assign n6091 = n492 & ~n6090;
  assign n6092 = n294 & ~n4023;
  assign n6093 = n408 & n6092;
  assign n6094 = ~n5824 & n6093;
  assign n6095 = ~n1325 & n5872;
  assign n6096 = n2623 & ~n6095;
  assign n6097 = ~n629 & ~n5027;
  assign n6098 = ~n4773 & n6097;
  assign n6099 = ~n6094 & n6098;
  assign n6100 = ~n1619 & n5486;
  assign n6101 = ~n6096 & n6100;
  assign n6102 = n6099 & n6101;
  assign n6103 = n851 & n4856;
  assign n6104 = n5871 & n6103;
  assign n6105 = ~n6091 & n6102;
  assign n6106 = n6104 & n6105;
  assign n6107 = n5189 & n6106;
  assign po058 = ~n5759 | ~n6107;
  assign n6109 = n533 & n5472;
  assign n6110 = n5232 & n6109;
  assign n6111 = n5451 & n6093;
  assign n6112 = n408 & n5474;
  assign n6113 = ~n6110 & ~n6112;
  assign n6114 = ~n2621 & n6113;
  assign n6115 = ~n6111 & n6114;
  assign n6116 = n4432 & n6115;
  assign n6117 = n2617 & n6116;
  assign n6118 = n5710 & n6117;
  assign po059 = ~n5610 | ~n6118;
  assign n6120 = ~n4047 & n5758;
  assign n6121 = n5949 & n6120;
  assign po060 = ~n5700 | ~n6121;
  assign n6123 = ~n2774 & n5257;
  assign n6124 = n4066 & n6123;
  assign n6125 = n1093 & ~n6124;
  assign n6126 = ~n4927 & ~n6125;
  assign n6127 = ~pi027 & ~n6126;
  assign n6128 = n5835 & n5836;
  assign n6129 = ~n4771 & ~n6128;
  assign n6130 = ~n3545 & n6129;
  assign n6131 = ~n1031 & n6130;
  assign n6132 = ~n1980 & n4919;
  assign n6133 = n6131 & n6132;
  assign n6134 = n5011 & n6133;
  assign n6135 = n5421 & n5762;
  assign n6136 = ~n5877 & n5978;
  assign n6137 = n6135 & n6136;
  assign n6138 = n6134 & n6137;
  assign po061 = n6127 | ~n6138;
  assign n6140 = pi027 & n2783;
  assign n6141 = n1338 & ~n5819;
  assign n6142 = ~n2590 & ~n3226;
  assign n6143 = ~n6141 & n6142;
  assign n6144 = n415 & n6143;
  assign n6145 = n3723 & n6144;
  assign n6146 = ~n6140 & n6145;
  assign po062 = ~n5808 | ~n6146;
  assign po063 = ~n3291 | n5436;
  assign n6149 = n487 & n668;
  assign n6150 = ~n2275 & ~n6149;
  assign n6151 = ~pi022 & ~n6150;
  assign n6152 = pi022 & n1857;
  assign n6153 = ~pi122 & ~n3037;
  assign n6154 = n2307 & n6153;
  assign n6155 = pi122 & n1078;
  assign n6156 = ~n357 & n6155;
  assign n6157 = n5382 & n6156;
  assign n6158 = ~n6154 & ~n6157;
  assign n6159 = pi122 & n386;
  assign n6160 = ~n1071 & ~n6159;
  assign n6161 = n1387 & ~n6160;
  assign n6162 = ~n973 & n1027;
  assign n6163 = ~n410 & ~n1071;
  assign n6164 = ~pi023 & ~n6163;
  assign n6165 = ~n568 & ~n575;
  assign n6166 = ~n6162 & n6165;
  assign n6167 = ~n6164 & n6166;
  assign n6168 = n362 & ~n6167;
  assign n6169 = ~n3080 & ~n3276;
  assign n6170 = ~n6168 & n6169;
  assign n6171 = ~n885 & ~n3090;
  assign n6172 = n6170 & n6171;
  assign n6173 = n5553 & ~n6152;
  assign n6174 = ~n6161 & n6173;
  assign n6175 = ~n1903 & n6172;
  assign n6176 = n6174 & n6175;
  assign n6177 = ~n6151 & n6176;
  assign n6178 = ~n6158 & n6177;
  assign n6179 = n293 & ~n6178;
  assign n6180 = n507 & n1500;
  assign n6181 = ~n1930 & n2770;
  assign n6182 = n4426 & n4808;
  assign n6183 = ~n6180 & n6182;
  assign n6184 = n6181 & n6183;
  assign n6185 = n5691 & n6184;
  assign n6186 = n492 & ~n6185;
  assign n6187 = n315 & n476;
  assign n6188 = n3055 & ~n3060;
  assign n6189 = n484 & n1387;
  assign n6190 = ~n2242 & ~n6189;
  assign n6191 = ~pi122 & ~n6190;
  assign n6192 = ~n990 & n1521;
  assign n6193 = n336 & n781;
  assign n6194 = ~n1571 & ~n6193;
  assign n6195 = n1228 & ~n6194;
  assign n6196 = n317 & n455;
  assign n6197 = ~n6195 & ~n6196;
  assign n6198 = ~pi044 & n391;
  assign n6199 = n603 & ~n1848;
  assign n6200 = ~pi065 & n3062;
  assign n6201 = ~pi020 & n3045;
  assign n6202 = ~n5579 & ~n6201;
  assign n6203 = n349 & n528;
  assign n6204 = ~n799 & n1435;
  assign n6205 = ~n1103 & ~n2656;
  assign n6206 = ~n6204 & n6205;
  assign n6207 = pi122 & ~n6206;
  assign n6208 = n476 & n2097;
  assign n6209 = pi022 & ~pi044;
  assign n6210 = ~n381 & ~n6209;
  assign n6211 = n417 & n6210;
  assign n6212 = n1387 & n6211;
  assign n6213 = ~n5559 & ~n6212;
  assign n6214 = n293 & ~n6213;
  assign n6215 = ~pi044 & pi122;
  assign n6216 = n484 & n6215;
  assign n6217 = n355 & n6216;
  assign n6218 = ~n6208 & ~n6217;
  assign n6219 = ~n6214 & n6218;
  assign n6220 = ~n6187 & ~n6203;
  assign n6221 = ~n1268 & n6220;
  assign n6222 = ~n1271 & ~n3319;
  assign n6223 = n6221 & n6222;
  assign n6224 = ~n6198 & n6223;
  assign n6225 = n6202 & n6224;
  assign n6226 = ~n1505 & n3904;
  assign n6227 = ~n6192 & n6197;
  assign n6228 = ~n6199 & ~n6200;
  assign n6229 = n6227 & n6228;
  assign n6230 = n6225 & n6226;
  assign n6231 = n2372 & ~n3056;
  assign n6232 = ~n6188 & ~n6191;
  assign n6233 = n6231 & n6232;
  assign n6234 = n6229 & n6230;
  assign n6235 = n5682 & ~n6207;
  assign n6236 = n6219 & n6235;
  assign n6237 = n6233 & n6234;
  assign n6238 = n6236 & n6237;
  assign n6239 = ~n6179 & n6238;
  assign n6240 = ~n6186 & n6239;
  assign n6241 = ~pi045 & ~n6240;
  assign n6242 = n1029 & n2646;
  assign n6243 = n5452 & n5816;
  assign n6244 = n1783 & n5457;
  assign n6245 = ~n5456 & ~n6244;
  assign n6246 = n6243 & ~n6245;
  assign n6247 = n454 & n5831;
  assign n6248 = ~n6246 & ~n6247;
  assign n6249 = ~n5814 & n6248;
  assign n6250 = ~n2357 & ~n2669;
  assign n6251 = ~n807 & ~n1463;
  assign n6252 = ~n2388 & n6251;
  assign n6253 = ~n2880 & n6252;
  assign n6254 = n6250 & n6253;
  assign n6255 = ~pi045 & ~n6254;
  assign n6256 = n4207 & n6249;
  assign n6257 = n3374 & n6256;
  assign n6258 = ~n6255 & n6257;
  assign n6259 = n330 & ~n6258;
  assign n6260 = n1673 & ~n5850;
  assign n6261 = n1132 & n4427;
  assign n6262 = ~n2094 & ~n6261;
  assign n6263 = n4414 & n6262;
  assign n6264 = ~n6260 & n6263;
  assign n6265 = n302 & n3368;
  assign n6266 = n6264 & ~n6265;
  assign n6267 = n1668 & ~n4095;
  assign n6268 = n628 & n789;
  assign n6269 = n368 & n467;
  assign n6270 = ~n441 & ~n6269;
  assign n6271 = n1064 & n1638;
  assign n6272 = n599 & n3757;
  assign n6273 = n566 & n6272;
  assign n6274 = ~n2698 & ~n6273;
  assign n6275 = ~pi039 & ~n6274;
  assign n6276 = ~n6271 & ~n6275;
  assign n6277 = n775 & n1228;
  assign n6278 = ~n3262 & ~n6277;
  assign n6279 = ~pi045 & ~n6278;
  assign n6280 = ~n1499 & ~n6268;
  assign n6281 = n6270 & n6280;
  assign n6282 = n6276 & ~n6279;
  assign n6283 = n6281 & n6282;
  assign n6284 = ~n3818 & ~n6267;
  assign n6285 = n6283 & n6284;
  assign n6286 = ~pi006 & ~n687;
  assign n6287 = n5831 & ~n6286;
  assign n6288 = ~n5443 & n5471;
  assign n6289 = n5815 & ~n6288;
  assign n6290 = ~n6287 & ~n6289;
  assign n6291 = n2646 & ~n6290;
  assign n6292 = ~pi045 & ~n5447;
  assign n6293 = ~n5462 & ~n6292;
  assign n6294 = n572 & n5817;
  assign n6295 = ~n6293 & n6294;
  assign n6296 = ~n6291 & ~n6295;
  assign n6297 = pi029 & ~n6296;
  assign n6298 = n533 & n1228;
  assign n6299 = ~pi011 & ~n302;
  assign n6300 = n5455 & n6299;
  assign n6301 = n4029 & ~n6244;
  assign n6302 = ~n6300 & n6301;
  assign n6303 = ~n350 & ~n6302;
  assign n6304 = n5816 & ~n6303;
  assign n6305 = pi029 & n2646;
  assign n6306 = n293 & n6305;
  assign n6307 = n6304 & n6306;
  assign n6308 = ~n6298 & ~n6307;
  assign n6309 = ~n6297 & n6308;
  assign n6310 = ~n5757 & n6309;
  assign n6311 = n4404 & n6310;
  assign n6312 = pi029 & n2682;
  assign n6313 = ~n1440 & n1952;
  assign n6314 = n5707 & ~n6313;
  assign n6315 = n740 & n3784;
  assign n6316 = ~pi045 & n593;
  assign n6317 = n568 & n6316;
  assign n6318 = pi013 & n1008;
  assign n6319 = ~pi011 & n6318;
  assign n6320 = n2646 & n5661;
  assign n6321 = n311 & n5604;
  assign n6322 = n1357 & n6321;
  assign n6323 = ~n511 & ~n933;
  assign n6324 = n354 & n4405;
  assign n6325 = ~n6323 & n6324;
  assign n6326 = ~n2580 & ~n3736;
  assign n6327 = ~n1798 & n6326;
  assign n6328 = n408 & ~n6327;
  assign n6329 = n1694 & ~n4088;
  assign n6330 = ~n1777 & n2584;
  assign n6331 = ~pi056 & n5703;
  assign n6332 = pi044 & n4385;
  assign n6333 = ~n391 & ~n1901;
  assign n6334 = n6332 & ~n6333;
  assign n6335 = ~n1584 & ~n6322;
  assign n6336 = ~n3859 & ~n3887;
  assign n6337 = ~n6320 & n6336;
  assign n6338 = ~n6319 & n6335;
  assign n6339 = ~n6325 & n6338;
  assign n6340 = n3908 & n6337;
  assign n6341 = ~n5702 & ~n6317;
  assign n6342 = ~n6330 & ~n6331;
  assign n6343 = n6341 & n6342;
  assign n6344 = n6339 & n6340;
  assign n6345 = ~n5385 & ~n6242;
  assign n6346 = ~n6329 & ~n6334;
  assign n6347 = n6345 & n6346;
  assign n6348 = n6343 & n6344;
  assign n6349 = ~n2369 & n3271;
  assign n6350 = ~n6312 & ~n6314;
  assign n6351 = ~n6315 & n6350;
  assign n6352 = n6348 & n6349;
  assign n6353 = ~n6328 & n6347;
  assign n6354 = n6352 & n6353;
  assign n6355 = n6311 & n6351;
  assign n6356 = n6354 & n6355;
  assign n6357 = n6285 & n6356;
  assign n6358 = ~n6259 & n6266;
  assign n6359 = n6357 & n6358;
  assign n6360 = ~n4424 & n6359;
  assign po065 = n6241 | ~n6360;
  assign n6362 = ~n2504 & ~n3225;
  assign n6363 = ~n2178 & n6362;
  assign n6364 = n6035 & n6363;
  assign n6365 = ~n2844 & n6364;
  assign n6366 = n2930 & n6365;
  assign n6367 = n3047 & n5520;
  assign n6368 = n2786 & n6367;
  assign n6369 = n2248 & n6368;
  assign n6370 = n2259 & ~n5560;
  assign n6371 = n5557 & n6370;
  assign n6372 = n293 & ~n6371;
  assign n6373 = ~n1420 & ~n2180;
  assign n6374 = ~n2898 & n6373;
  assign n6375 = n6197 & n6374;
  assign n6376 = n6366 & n6375;
  assign n6377 = n6369 & n6376;
  assign n6378 = ~n6372 & n6377;
  assign n6379 = ~pi045 & ~n6378;
  assign n6380 = n5497 & n6250;
  assign n6381 = n318 & n1598;
  assign n6382 = n2193 & ~n6381;
  assign n6383 = n6380 & n6382;
  assign n6384 = n6305 & ~n6383;
  assign n6385 = ~pi023 & n420;
  assign n6386 = ~n486 & ~n6385;
  assign n6387 = n3642 & ~n6386;
  assign n6388 = ~n1875 & ~n6387;
  assign n6389 = pi018 & ~n6388;
  assign n6390 = ~n799 & n1092;
  assign n6391 = n1070 & n6316;
  assign n6392 = pi122 & n4405;
  assign n6393 = n3621 & n6392;
  assign n6394 = ~n6391 & ~n6393;
  assign n6395 = ~pi021 & ~n6394;
  assign n6396 = n1388 & n4396;
  assign n6397 = ~n1044 & ~n6396;
  assign n6398 = ~pi045 & ~n990;
  assign n6399 = ~n1952 & n6398;
  assign n6400 = ~n1952 & n5707;
  assign n6401 = n492 & n811;
  assign n6402 = n2774 & n6401;
  assign n6403 = pi022 & n812;
  assign n6404 = n411 & n2381;
  assign n6405 = ~pi045 & n480;
  assign n6406 = n732 & n6405;
  assign n6407 = ~n492 & ~n6305;
  assign n6408 = n797 & ~n6407;
  assign n6409 = n376 & n555;
  assign n6410 = ~n6406 & ~n6409;
  assign n6411 = ~n6402 & n6410;
  assign n6412 = ~n6408 & n6411;
  assign n6413 = ~n6318 & ~n6404;
  assign n6414 = n6412 & n6413;
  assign n6415 = ~n709 & n6414;
  assign n6416 = ~n2721 & n6415;
  assign n6417 = ~n6390 & n6397;
  assign n6418 = ~n6399 & ~n6400;
  assign n6419 = ~n6403 & n6418;
  assign n6420 = n6416 & n6417;
  assign n6421 = ~n5761 & ~n6389;
  assign n6422 = ~n6395 & n6421;
  assign n6423 = n6419 & n6420;
  assign n6424 = ~n3623 & n4054;
  assign n6425 = n6423 & n6424;
  assign n6426 = n2384 & n6422;
  assign n6427 = ~n6384 & n6426;
  assign n6428 = n6425 & n6427;
  assign n6429 = ~n6379 & n6428;
  assign n6430 = n5713 & n6429;
  assign n6431 = ~n2388 & ~n2539;
  assign n6432 = n6305 & ~n6431;
  assign n6433 = n349 & n6332;
  assign n6434 = n2326 & n6433;
  assign n6435 = ~n667 & ~n2230;
  assign n6436 = n2228 & ~n6435;
  assign n6437 = n2233 & ~n6436;
  assign n6438 = ~n2979 & ~n3728;
  assign n6439 = ~n6437 & n6438;
  assign n6440 = ~pi045 & ~n6439;
  assign n6441 = ~n1900 & ~n3460;
  assign n6442 = ~pi044 & ~n6441;
  assign n6443 = ~n375 & ~n550;
  assign n6444 = n377 & ~n6443;
  assign n6445 = ~n6442 & ~n6444;
  assign n6446 = n4385 & ~n6445;
  assign n6447 = n476 & n6332;
  assign n6448 = n479 & n6447;
  assign n6449 = ~pi045 & n2233;
  assign n6450 = n1418 & n6449;
  assign n6451 = ~n6434 & ~n6448;
  assign n6452 = ~n6450 & n6451;
  assign n6453 = ~n6446 & n6452;
  assign n6454 = ~n6440 & n6453;
  assign n6455 = ~pi122 & ~n5783;
  assign n6456 = n4000 & ~n6455;
  assign n6457 = n349 & ~n6456;
  assign n6458 = ~pi044 & ~n2876;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = ~n3077 & n6459;
  assign n6461 = ~n3041 & n6460;
  assign n6462 = n6219 & n6461;
  assign n6463 = ~pi045 & ~n6462;
  assign n6464 = n2784 & ~n5633;
  assign n6465 = n811 & ~n6464;
  assign n6466 = ~n2936 & ~n5558;
  assign n6467 = n4405 & ~n6466;
  assign n6468 = n310 & n5604;
  assign n6469 = n2290 & n4385;
  assign n6470 = ~n6468 & ~n6469;
  assign n6471 = n416 & ~n6470;
  assign n6472 = ~n2942 & n6392;
  assign n6473 = ~n1598 & ~n2010;
  assign n6474 = n4385 & ~n6473;
  assign n6475 = n811 & n957;
  assign n6476 = n310 & n6475;
  assign n6477 = ~n6474 & ~n6476;
  assign n6478 = n475 & ~n6477;
  assign n6479 = ~n6471 & ~n6478;
  assign n6480 = ~n6432 & n6479;
  assign n6481 = ~n6467 & n6480;
  assign n6482 = ~n6465 & ~n6472;
  assign n6483 = n6481 & n6482;
  assign n6484 = n6454 & n6483;
  assign n6485 = ~n6463 & n6484;
  assign n6486 = ~n2291 & n6333;
  assign n6487 = n6332 & ~n6486;
  assign n6488 = ~pi045 & ~n6215;
  assign n6489 = n2873 & n6488;
  assign n6490 = ~n6487 & ~n6489;
  assign n6491 = n6485 & n6490;
  assign n6492 = ~n2583 & ~n6330;
  assign n6493 = n567 & n5491;
  assign n6494 = n1246 & ~n3088;
  assign n6495 = n372 & ~n2284;
  assign n6496 = ~pi029 & n3826;
  assign n6497 = ~n6494 & ~n6495;
  assign n6498 = ~n3808 & n6497;
  assign n6499 = ~n6496 & n6498;
  assign n6500 = pi122 & ~n6499;
  assign n6501 = ~n990 & n3637;
  assign n6502 = ~pi023 & ~n1427;
  assign n6503 = n949 & ~n2252;
  assign n6504 = ~n6502 & ~n6503;
  assign n6505 = n416 & ~n6504;
  assign n6506 = n3891 & n5494;
  assign n6507 = n2311 & ~n6506;
  assign n6508 = ~n6501 & n6507;
  assign n6509 = ~n6505 & n6508;
  assign n6510 = ~n6500 & n6509;
  assign n6511 = ~pi045 & ~n6510;
  assign n6512 = n827 & n4385;
  assign n6513 = ~n835 & n6512;
  assign n6514 = ~n2589 & ~n5233;
  assign n6515 = n1190 & n1531;
  assign n6516 = n492 & n6515;
  assign n6517 = n1294 & n6516;
  assign n6518 = n6514 & ~n6517;
  assign n6519 = ~n6513 & n6518;
  assign n6520 = ~n5489 & n6519;
  assign n6521 = ~n6493 & n6520;
  assign n6522 = n6492 & n6521;
  assign n6523 = ~n6511 & n6522;
  assign n6524 = n1337 & n6247;
  assign n6525 = n5819 & ~n6246;
  assign n6526 = ~n5492 & n6525;
  assign n6527 = n492 & ~n6526;
  assign n6528 = n5452 & n6092;
  assign n6529 = n5437 & ~n5466;
  assign n6530 = ~n533 & ~n5470;
  assign n6531 = ~n6529 & n6530;
  assign n6532 = pi029 & ~n6531;
  assign n6533 = ~n6528 & ~n6532;
  assign n6534 = n537 & ~n6533;
  assign n6535 = n293 & n4427;
  assign n6536 = n6304 & n6535;
  assign n6537 = ~n6524 & ~n6536;
  assign n6538 = ~n6534 & n6537;
  assign n6539 = ~n6527 & n6538;
  assign n6540 = n6523 & n6539;
  assign n6541 = n585 & n2487;
  assign n6542 = n1833 & ~n6541;
  assign n6543 = n329 & ~n6542;
  assign n6544 = n1241 & ~n6386;
  assign n6545 = ~n3251 & ~n6544;
  assign n6546 = n1624 & ~n6545;
  assign n6547 = n1590 & n1682;
  assign n6548 = n949 & n1260;
  assign n6549 = ~n937 & ~n6547;
  assign n6550 = ~n3640 & n6549;
  assign n6551 = ~n6548 & n6550;
  assign n6552 = ~n2275 & n6551;
  assign n6553 = n315 & ~n6552;
  assign n6554 = ~n4452 & ~n6329;
  assign n6555 = n2567 & ~n4169;
  assign n6556 = n1338 & ~n6555;
  assign n6557 = n6554 & ~n6556;
  assign n6558 = ~n1865 & n4180;
  assign n6559 = ~n6546 & n6558;
  assign n6560 = ~n6553 & n6559;
  assign n6561 = n6557 & n6560;
  assign n6562 = n1228 & n1699;
  assign n6563 = ~n1789 & ~n6562;
  assign n6564 = n692 & ~n6563;
  assign n6565 = n693 & n4074;
  assign n6566 = pi011 & ~n2487;
  assign n6567 = n1667 & ~n2488;
  assign n6568 = ~n6566 & n6567;
  assign n6569 = ~n705 & n2543;
  assign n6570 = ~n448 & ~n1702;
  assign n6571 = n1704 & ~n6570;
  assign n6572 = n329 & n4094;
  assign n6573 = ~n1694 & ~n6572;
  assign n6574 = n585 & ~n6573;
  assign n6575 = ~n3312 & ~n3530;
  assign n6576 = ~n4152 & n6575;
  assign n6577 = n1754 & ~n6576;
  assign n6578 = ~n1720 & ~n6571;
  assign n6579 = ~n2535 & ~n6569;
  assign n6580 = n6578 & n6579;
  assign n6581 = ~n1707 & ~n2595;
  assign n6582 = ~n3573 & ~n6565;
  assign n6583 = ~n6568 & n6582;
  assign n6584 = n6580 & n6581;
  assign n6585 = n4839 & ~n6564;
  assign n6586 = ~n6577 & n6585;
  assign n6587 = n6583 & n6584;
  assign n6588 = ~n6574 & n6587;
  assign n6589 = n3523 & n6586;
  assign n6590 = n6588 & n6589;
  assign n6591 = n2626 & n6590;
  assign n6592 = ~n6543 & n6561;
  assign n6593 = n6591 & n6592;
  assign n6594 = n5448 & n5816;
  assign n6595 = n5677 & n6594;
  assign n6596 = ~n1583 & ~n2880;
  assign n6597 = n1002 & n6596;
  assign n6598 = n740 & ~n6597;
  assign n6599 = n415 & ~n6598;
  assign n6600 = n1673 & ~n4924;
  assign n6601 = ~pi027 & n5899;
  assign n6602 = n1264 & n1480;
  assign n6603 = ~n6600 & ~n6602;
  assign n6604 = ~n6601 & n6603;
  assign n6605 = ~n6312 & n6604;
  assign n6606 = n6599 & n6605;
  assign n6607 = n403 & n1396;
  assign n6608 = ~n640 & ~n6607;
  assign n6609 = n6206 & n6608;
  assign n6610 = n2653 & n6609;
  assign n6611 = n4385 & ~n6610;
  assign n6612 = ~pi044 & n406;
  assign n6613 = ~n2793 & ~n6612;
  assign n6614 = n3273 & ~n5495;
  assign n6615 = n6613 & n6614;
  assign n6616 = n6290 & n6615;
  assign n6617 = n2772 & n6616;
  assign n6618 = n4427 & ~n6617;
  assign n6619 = ~n468 & n4205;
  assign n6620 = n330 & ~n6619;
  assign n6621 = ~n621 & ~n4796;
  assign n6622 = n1718 & ~n6621;
  assign n6623 = n479 & n751;
  assign n6624 = pi122 & n4427;
  assign n6625 = n6623 & n6624;
  assign n6626 = n1728 & ~n1746;
  assign n6627 = ~n4563 & ~n6626;
  assign n6628 = n4059 & ~n6627;
  assign n6629 = ~n4073 & ~n6625;
  assign n6630 = ~n6595 & n6629;
  assign n6631 = ~n5368 & n6630;
  assign n6632 = ~n6628 & n6631;
  assign n6633 = ~n6622 & n6632;
  assign n6634 = ~n6620 & n6633;
  assign n6635 = n5760 & ~n6618;
  assign n6636 = n6634 & n6635;
  assign n6637 = n6606 & ~n6611;
  assign n6638 = n6636 & n6637;
  assign n6639 = n6285 & n6638;
  assign n6640 = n6593 & n6639;
  assign n6641 = n6491 & n6640;
  assign n6642 = n6540 & n6641;
  assign po066 = ~n6430 | ~n6642;
  assign n6644 = n699 & n6316;
  assign n6645 = n492 & n1225;
  assign n6646 = n4422 & ~n6645;
  assign n6647 = n4388 & ~n6646;
  assign n6648 = n2381 & ~n2836;
  assign n6649 = n1539 & n6648;
  assign n6650 = n743 & ~n6215;
  assign n6651 = n329 & n6650;
  assign n6652 = n403 & n6651;
  assign n6653 = ~n2764 & ~n6652;
  assign n6654 = n2365 & ~n6653;
  assign n6655 = ~n6649 & ~n6654;
  assign n6656 = n4403 & n6655;
  assign n6657 = ~n6647 & n6656;
  assign n6658 = n1076 & n1516;
  assign n6659 = ~n937 & ~n2848;
  assign n6660 = n2271 & n6659;
  assign n6661 = ~n2932 & n6660;
  assign n6662 = n416 & ~n6661;
  assign n6663 = ~n878 & n6608;
  assign n6664 = n2654 & n6663;
  assign n6665 = pi122 & ~n6664;
  assign n6666 = n2720 & n3103;
  assign n6667 = n2565 & ~n3060;
  assign n6668 = n507 & n2092;
  assign n6669 = ~n6667 & ~n6668;
  assign n6670 = pi022 & ~n6669;
  assign n6671 = pi065 & n3062;
  assign n6672 = ~pi044 & ~n2875;
  assign n6673 = n333 & n335;
  assign n6674 = n480 & n6673;
  assign n6675 = n350 & n2000;
  assign n6676 = n375 & ~n2294;
  assign n6677 = ~n2001 & ~n6676;
  assign n6678 = n306 & ~n6677;
  assign n6679 = ~n1431 & ~n6675;
  assign n6680 = ~n6674 & n6679;
  assign n6681 = ~n3058 & n6680;
  assign n6682 = ~n1972 & ~n6678;
  assign n6683 = n6681 & n6682;
  assign n6684 = ~n1506 & ~n6672;
  assign n6685 = n6683 & n6684;
  assign n6686 = ~n1726 & ~n2988;
  assign n6687 = n5520 & ~n6658;
  assign n6688 = n6686 & n6687;
  assign n6689 = ~n6666 & n6685;
  assign n6690 = ~n6671 & n6689;
  assign n6691 = n2378 & n6688;
  assign n6692 = n6690 & n6691;
  assign n6693 = ~n2236 & n5657;
  assign n6694 = ~n6670 & n6693;
  assign n6695 = ~n6665 & n6692;
  assign n6696 = n6694 & n6695;
  assign n6697 = n6366 & ~n6662;
  assign n6698 = n6696 & n6697;
  assign n6699 = ~pi045 & ~n6698;
  assign n6700 = n330 & ~n1833;
  assign n6701 = n2646 & ~n3028;
  assign n6702 = n492 & ~n3100;
  assign n6703 = n5704 & ~n6702;
  assign n6704 = ~pi056 & ~n6703;
  assign n6705 = ~n1513 & n3110;
  assign n6706 = ~n1294 & ~n1328;
  assign n6707 = n6616 & n6706;
  assign n6708 = n6705 & n6707;
  assign n6709 = n4427 & ~n6708;
  assign n6710 = n349 & ~n3457;
  assign n6711 = ~n1900 & n2324;
  assign n6712 = ~n6710 & n6711;
  assign n6713 = n811 & ~n6712;
  assign n6714 = pi023 & pi122;
  assign n6715 = n5547 & ~n6714;
  assign n6716 = ~n2845 & ~n4592;
  assign n6717 = n1243 & ~n6716;
  assign n6718 = ~n1261 & ~n6717;
  assign n6719 = ~n6715 & n6718;
  assign n6720 = n4405 & ~n6719;
  assign n6721 = ~n1919 & ~n5594;
  assign n6722 = n1571 & n6721;
  assign n6723 = ~n752 & ~n6722;
  assign n6724 = n6624 & ~n6723;
  assign n6725 = n602 & ~n6594;
  assign n6726 = ~n1886 & n6725;
  assign n6727 = n5677 & ~n6726;
  assign n6728 = ~n797 & ~n6381;
  assign n6729 = ~n1309 & n6728;
  assign n6730 = ~n1464 & n6729;
  assign n6731 = ~n1501 & n1627;
  assign n6732 = n6730 & n6731;
  assign n6733 = n6305 & ~n6732;
  assign n6734 = n853 & n1668;
  assign n6735 = n1915 & n6398;
  assign n6736 = n2291 & n6332;
  assign n6737 = n419 & n2381;
  assign n6738 = n972 & n6737;
  assign n6739 = n1074 & n5412;
  assign n6740 = n362 & n6739;
  assign n6741 = ~n6738 & ~n6740;
  assign n6742 = ~pi019 & ~n6741;
  assign n6743 = ~n6724 & ~n6736;
  assign n6744 = ~n6734 & ~n6735;
  assign n6745 = n6743 & n6744;
  assign n6746 = ~n2382 & ~n3364;
  assign n6747 = ~n6713 & n6746;
  assign n6748 = ~n6644 & n6745;
  assign n6749 = ~n6742 & n6748;
  assign n6750 = ~n3857 & n6747;
  assign n6751 = n6749 & n6750;
  assign n6752 = n6554 & ~n6720;
  assign n6753 = ~n6727 & ~n6733;
  assign n6754 = n6752 & n6753;
  assign n6755 = ~n6704 & n6751;
  assign n6756 = n6754 & n6755;
  assign n6757 = ~n6700 & ~n6709;
  assign n6758 = n6756 & n6757;
  assign n6759 = n5675 & n6454;
  assign n6760 = n6758 & n6759;
  assign n6761 = n6266 & ~n6701;
  assign n6762 = n6760 & n6761;
  assign n6763 = ~n6699 & n6762;
  assign n6764 = n6540 & n6657;
  assign po067 = ~n6763 | ~n6764;
  assign n6766 = pi029 & n472;
  assign n6767 = n6606 & ~n6766;
  assign n6768 = n330 & ~n4205;
  assign n6769 = n4058 & n6562;
  assign n6770 = n809 & n1241;
  assign n6771 = ~pi015 & n2575;
  assign n6772 = ~n1702 & ~n4563;
  assign n6773 = n4059 & ~n6772;
  assign n6774 = ~n3636 & ~n6770;
  assign n6775 = ~n6267 & n6774;
  assign n6776 = ~n6769 & ~n6773;
  assign n6777 = n6775 & n6776;
  assign n6778 = ~n6768 & ~n6771;
  assign n6779 = n6777 & n6778;
  assign n6780 = n5986 & n6779;
  assign n6781 = ~n4043 & n6780;
  assign n6782 = n6492 & n6781;
  assign n6783 = n6767 & n6782;
  assign po068 = ~n6593 | ~n6783;
  assign n6785 = n1754 & ~n5176;
  assign n6786 = n1668 & ~n4096;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = ~n6700 & n6787;
  assign n6789 = n2587 & n6788;
  assign n6790 = n330 & ~n6249;
  assign n6791 = ~n3539 & ~n6790;
  assign n6792 = n3371 & n6791;
  assign n6793 = n6263 & n6792;
  assign n6794 = n6311 & n6557;
  assign n6795 = n6793 & n6794;
  assign n6796 = n6767 & n6795;
  assign n6797 = n6789 & n6796;
  assign po069 = ~n4429 | ~n6797;
  assign n6799 = n2654 & n6609;
  assign n6800 = n4385 & ~n6799;
  assign n6801 = n740 & n2880;
  assign n6802 = n329 & n5492;
  assign n6803 = ~pi029 & n6802;
  assign n6804 = n1724 & n4796;
  assign n6805 = ~n6623 & ~n6722;
  assign n6806 = n6624 & ~n6805;
  assign n6807 = n2773 & n6615;
  assign n6808 = n4427 & ~n6807;
  assign n6809 = ~n3532 & ~n5188;
  assign n6810 = pi029 & ~n6809;
  assign n6811 = ~n5027 & ~n6806;
  assign n6812 = ~n4060 & n6811;
  assign n6813 = ~n5374 & ~n6801;
  assign n6814 = ~n6804 & n6813;
  assign n6815 = ~n6771 & n6812;
  assign n6816 = ~n6785 & n6815;
  assign n6817 = ~n6487 & n6814;
  assign n6818 = n6816 & n6817;
  assign n6819 = ~n6808 & n6818;
  assign n6820 = n6283 & ~n6800;
  assign n6821 = ~n6803 & ~n6810;
  assign n6822 = n6820 & n6821;
  assign n6823 = n3376 & n6819;
  assign n6824 = n6264 & n6561;
  assign n6825 = n6823 & n6824;
  assign n6826 = n6822 & n6825;
  assign n6827 = n6485 & n6523;
  assign n6828 = n6826 & n6827;
  assign n6829 = n6657 & n6828;
  assign po070 = ~n6430 | ~n6829;
  assign n6831 = ~n470 & ~n5084;
  assign n6832 = n5819 & n6831;
  assign n6833 = ~n3538 & n6832;
  assign n6834 = n329 & ~n6833;
  assign n6835 = ~n574 & ~n6834;
  assign po071 = ~n6599 | ~n6835;
  assign n6837 = ~pi006 & pi029;
  assign n6838 = ~pi066 & n6837;
  assign n6839 = n782 & ~n6838;
  assign n6840 = n780 & ~n6839;
  assign n6841 = n329 & ~n6840;
  assign n6842 = n1029 & n1095;
  assign n6843 = n6276 & ~n6842;
  assign po073 = n6841 | ~n6843;
  assign n6845 = pi029 & ~n4207;
  assign n6846 = n6248 & ~n6845;
  assign n6847 = n329 & ~n6846;
  assign n6848 = ~n441 & ~n3369;
  assign n6849 = ~n5161 & n6848;
  assign n6850 = ~n6329 & n6849;
  assign n6851 = n6605 & n6850;
  assign n6852 = ~n6847 & n6851;
  assign po074 = ~n6789 | ~n6852;
  assign n6854 = ~n6243 & ~n6247;
  assign n6855 = n1338 & ~n6854;
  assign n6856 = ~n709 & ~n6269;
  assign po075 = n6855 | ~n6856;
  assign n6858 = ~n1760 & n2605;
  assign n6859 = pi029 & n3365;
  assign po076 = ~n6858 | n6859;
  assign n6861 = ~n1707 & ~n3673;
  assign n6862 = n330 & n3300;
  assign n6863 = n368 & n1705;
  assign n6864 = ~n3521 & ~n6863;
  assign n6865 = ~n2535 & ~n4231;
  assign n6866 = ~n2523 & n6865;
  assign n6867 = ~n2610 & ~n6862;
  assign n6868 = n6864 & n6867;
  assign n6869 = ~n2624 & n6866;
  assign n6870 = n6861 & n6869;
  assign n6871 = n6868 & n6870;
  assign po077 = ~n2493 | ~n6871;
  assign n6873 = n332 & n2543;
  assign n6874 = n6514 & ~n6873;
  assign n6875 = n3475 & n6874;
  assign n6876 = ~n6400 & n6875;
  assign po078 = ~n5710 | ~n6876;
  assign n6878 = n4590 & n5557;
  assign n6879 = n293 & ~n6878;
  assign n6880 = ~n5249 & n6369;
  assign n6881 = ~n1420 & ~n6879;
  assign n6882 = n6880 & n6881;
  assign n6883 = ~pi045 & ~n6882;
  assign n6884 = n1435 & n5503;
  assign n6885 = ~n6046 & ~n6607;
  assign n6886 = n2995 & n6885;
  assign n6887 = n4385 & ~n6886;
  assign n6888 = n4218 & n6613;
  assign n6889 = n4427 & ~n6888;
  assign n6890 = n802 & n2388;
  assign n6891 = pi028 & n6890;
  assign n6892 = pi039 & pi045;
  assign n6893 = n350 & n632;
  assign n6894 = n336 & n616;
  assign n6895 = ~pi005 & n6894;
  assign n6896 = n1392 & n6895;
  assign n6897 = ~n3484 & ~n6893;
  assign n6898 = ~n6896 & n6897;
  assign n6899 = ~pi122 & n6892;
  assign n6900 = ~n6898 & n6899;
  assign n6901 = n1952 & n5572;
  assign n6902 = n6398 & ~n6901;
  assign n6903 = ~n2952 & n4406;
  assign n6904 = n2095 & ~n6884;
  assign n6905 = ~n6891 & n6904;
  assign n6906 = n2722 & n6905;
  assign n6907 = ~n6900 & n6906;
  assign n6908 = ~n6902 & ~n6903;
  assign n6909 = n6907 & n6908;
  assign n6910 = ~n6887 & ~n6889;
  assign n6911 = n6909 & n6910;
  assign n6912 = n6491 & n6911;
  assign n6913 = n2857 & ~n4417;
  assign n6914 = n5596 & ~n6913;
  assign n6915 = n2863 & ~n6914;
  assign n6916 = ~n5597 & ~n6915;
  assign n6917 = n1134 & ~n5594;
  assign n6918 = ~n6332 & ~n6917;
  assign n6919 = ~n4418 & ~n6918;
  assign n6920 = n293 & n4394;
  assign n6921 = ~n2104 & ~n6920;
  assign n6922 = n5593 & ~n6921;
  assign n6923 = ~n1521 & ~n4425;
  assign n6924 = ~pi056 & ~n6923;
  assign n6925 = ~n1915 & ~n6924;
  assign n6926 = n492 & ~n6925;
  assign n6927 = ~n1227 & ~n1230;
  assign n6928 = ~n6922 & n6927;
  assign n6929 = ~n6919 & n6928;
  assign n6930 = ~n6926 & n6929;
  assign n6931 = n5608 & ~n6916;
  assign n6932 = n6930 & n6931;
  assign n6933 = ~pi021 & ~n642;
  assign n6934 = ~n431 & n566;
  assign n6935 = ~n3639 & n6934;
  assign n6936 = ~n6933 & n6935;
  assign n6937 = ~n669 & ~n6936;
  assign n6938 = n6737 & ~n6937;
  assign n6939 = n2043 & ~n6938;
  assign n6940 = n6932 & n6939;
  assign n6941 = n6912 & n6940;
  assign po081 = n6883 | ~n6941;
  assign n6943 = n5357 & ~n6319;
  assign po079 = po081 | ~n6943;
  assign n6945 = ~n302 & ~n3228;
  assign n6946 = n677 & n6945;
  assign n6947 = pi020 & po123;
  assign n6948 = n1338 & n3055;
  assign n6949 = ~pi019 & ~n6933;
  assign n6950 = pi018 & ~n3576;
  assign n6951 = ~n6949 & ~n6950;
  assign n6952 = pi020 & n315;
  assign n6953 = ~n6951 & n6952;
  assign n6954 = n390 & n6953;
  assign n6955 = ~n6948 & ~n6954;
  assign n6956 = n1721 & ~n6947;
  assign n6957 = ~n4047 & n6956;
  assign po082 = ~n6955 | ~n6957;
  assign n6959 = ~n1044 & ~n6946;
  assign po080 = po082 | ~n6959;
  assign po083 = po081 | n6948;
  assign n6962 = ~n2545 & ~n3081;
  assign n6963 = ~pi044 & ~n6962;
  assign n6964 = pi044 & n3267;
  assign n6965 = n1418 & n6964;
  assign n6966 = ~n6149 & ~n6965;
  assign n6967 = ~n6963 & n6966;
  assign n6968 = n2277 & n6967;
  assign n6969 = pi122 & ~n6968;
  assign n6970 = n5044 & n5552;
  assign n6971 = ~n6969 & n6970;
  assign n6972 = n293 & ~n6971;
  assign n6973 = n6880 & ~n6972;
  assign n6974 = ~pi045 & ~n6973;
  assign n6975 = n354 & n4592;
  assign n6976 = n3082 & ~n6975;
  assign n6977 = ~n5554 & n6976;
  assign n6978 = n4396 & ~n6977;
  assign n6979 = n933 & n6324;
  assign n6980 = n4406 & n5014;
  assign n6981 = ~pi044 & n4385;
  assign n6982 = n483 & n6981;
  assign n6983 = ~n6980 & ~n6982;
  assign n6984 = pi019 & ~n6983;
  assign n6985 = n1419 & n6984;
  assign n6986 = pi019 & pi122;
  assign n6987 = ~pi045 & ~n6986;
  assign n6988 = n1420 & n6987;
  assign n6989 = ~n6946 & ~n6979;
  assign n6990 = ~n6985 & n6989;
  assign n6991 = ~n6988 & n6990;
  assign n6992 = n6397 & n6991;
  assign n6993 = n6955 & ~n6978;
  assign n6994 = n6992 & n6993;
  assign n6995 = ~n6974 & n6994;
  assign po084 = ~n6941 | ~n6995;
  assign po086 = n2094 | ~n6932;
  assign n6998 = ~pi013 & ~n589;
  assign n6999 = n320 & ~n6998;
  assign n7000 = ~pi022 & n1723;
  assign n7001 = ~n528 & ~n2000;
  assign n7002 = ~pi006 & n551;
  assign n7003 = ~n7001 & n7002;
  assign n7004 = ~n6999 & ~n7003;
  assign n7005 = ~n3250 & n7004;
  assign n7006 = ~n3320 & n7005;
  assign n7007 = ~n3746 & ~n7000;
  assign n7008 = n7006 & n7007;
  assign n7009 = n1974 & ~n4251;
  assign n7010 = n7008 & n7009;
  assign n7011 = n2410 & n7010;
  assign n7012 = n1946 & ~n4249;
  assign po087 = ~n7011 | ~n7012;
  assign n7014 = ~n802 & n4537;
  assign n7015 = n1316 & ~n7014;
  assign n7016 = ~n1269 & ~n2917;
  assign n7017 = ~n1231 & n7016;
  assign n7018 = n1497 & n7017;
  assign n7019 = ~n7015 & n7018;
  assign n7020 = n3030 & n7019;
  assign n7021 = n1302 & n1306;
  assign n7022 = ~n1535 & ~n7021;
  assign n7023 = n1228 & n2724;
  assign n7024 = n791 & n1328;
  assign n7025 = ~n1377 & n1501;
  assign n7026 = ~n7024 & ~n7025;
  assign n7027 = ~n7023 & n7026;
  assign n7028 = ~n1528 & n4431;
  assign n7029 = n1376 & ~n1469;
  assign n7030 = n1326 & n2763;
  assign n7031 = n604 & ~n2827;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = n1167 & ~n1897;
  assign n7034 = n1243 & n3995;
  assign n7035 = ~n5669 & ~n7034;
  assign n7036 = ~n360 & ~n7035;
  assign n7037 = n1513 & n2677;
  assign n7038 = n791 & n1345;
  assign n7039 = ~n1187 & ~n7037;
  assign n7040 = n2608 & n7039;
  assign n7041 = ~n7038 & n7040;
  assign n7042 = ~n7036 & n7041;
  assign n7043 = n2312 & n2410;
  assign n7044 = n4617 & n7033;
  assign n7045 = n7043 & n7044;
  assign n7046 = n7028 & n7042;
  assign n7047 = ~n7029 & n7032;
  assign n7048 = n7046 & n7047;
  assign n7049 = n1156 & n7045;
  assign n7050 = ~n2469 & n7027;
  assign n7051 = n7049 & n7050;
  assign n7052 = n1458 & n7048;
  assign n7053 = n2869 & n3318;
  assign n7054 = n7022 & n7053;
  assign n7055 = n7051 & n7052;
  assign n7056 = n1349 & n7055;
  assign n7057 = n1415 & n7054;
  assign n7058 = n7056 & n7057;
  assign po088 = ~n7020 | ~n7058;
  assign n7060 = n2907 & n4162;
  assign n7061 = n3087 & ~n3090;
  assign n7062 = n293 & ~n7061;
  assign n7063 = n3059 & ~n7062;
  assign n7064 = ~n360 & ~n7063;
  assign n7065 = n329 & ~n3707;
  assign n7066 = ~n2302 & n2304;
  assign n7067 = n5944 & n7066;
  assign n7068 = n345 & ~n7067;
  assign n7069 = ~n1132 & ~n3872;
  assign n7070 = n492 & ~n7069;
  assign n7071 = ~pi023 & ~n3069;
  assign n7072 = n949 & n7071;
  assign n7073 = ~n1490 & ~n7072;
  assign n7074 = n938 & ~n7073;
  assign n7075 = ~n360 & n2717;
  assign n7076 = ~n1518 & n2720;
  assign n7077 = ~pi039 & n4385;
  assign n7078 = n2994 & n7077;
  assign n7079 = ~n1038 & ~n2958;
  assign n7080 = ~n1084 & n7079;
  assign n7081 = ~n1231 & ~n2993;
  assign n7082 = n7080 & n7081;
  assign n7083 = ~n1970 & ~n7070;
  assign n7084 = n7082 & n7083;
  assign n7085 = ~n887 & ~n3633;
  assign n7086 = n3977 & ~n5162;
  assign n7087 = ~n7074 & ~n7076;
  assign n7088 = ~n7078 & n7087;
  assign n7089 = n7085 & n7086;
  assign n7090 = n2964 & n7084;
  assign n7091 = n4174 & ~n7075;
  assign n7092 = n7090 & n7091;
  assign n7093 = n7088 & n7089;
  assign n7094 = ~n3041 & n7028;
  assign n7095 = n7093 & n7094;
  assign n7096 = ~n7065 & n7092;
  assign n7097 = ~n7068 & n7096;
  assign n7098 = n2956 & n7095;
  assign n7099 = n7097 & n7098;
  assign n7100 = n4226 & n7060;
  assign n7101 = ~n7064 & n7100;
  assign n7102 = n7099 & n7101;
  assign n7103 = n4297 & n7102;
  assign po089 = ~n2892 | ~n7103;
  assign n7105 = n630 & n1579;
  assign n7106 = ~pi031 & pi032;
  assign n7107 = ~n2701 & n7106;
  assign n7108 = ~n534 & n1095;
  assign n7109 = ~pi122 & n1883;
  assign n7110 = ~n1444 & ~n3058;
  assign n7111 = ~n360 & ~n7110;
  assign n7112 = n2928 & ~n7111;
  assign n7113 = ~n2185 & ~n7109;
  assign po100 = ~n7112 | ~n7113;
  assign n7115 = ~n2811 & ~n7108;
  assign n7116 = ~n7107 & n7115;
  assign po091 = po100 | ~n7116;
  assign po090 = n7105 | po091;
  assign n7119 = pi031 & ~n2701;
  assign n7120 = ~n534 & n740;
  assign n7121 = ~n2813 & ~n7120;
  assign po092 = n7119 | ~n7121;
  assign n7123 = ~n1571 & n3113;
  assign n7124 = n492 & ~n7123;
  assign n7125 = ~n1893 & n2861;
  assign n7126 = ~n6645 & n7125;
  assign n7127 = ~n4412 & n7126;
  assign n7128 = n4421 & n7127;
  assign n7129 = ~n1153 & ~n2036;
  assign n7130 = ~n5701 & n7129;
  assign n7131 = n5705 & n7130;
  assign n7132 = ~n7124 & n7131;
  assign n7133 = n7128 & n7132;
  assign n7134 = n1135 & ~n7133;
  assign n7135 = pi044 & n6624;
  assign n7136 = n376 & n7135;
  assign n7137 = n1171 & n7136;
  assign n7138 = n345 & n1190;
  assign n7139 = ~pi065 & n6332;
  assign n7140 = ~n7138 & ~n7139;
  assign n7141 = n2916 & ~n7140;
  assign n7142 = n518 & n6332;
  assign n7143 = n771 & n7142;
  assign n7144 = ~n7136 & ~n7143;
  assign n7145 = n1177 & ~n7144;
  assign n7146 = n492 & n1135;
  assign n7147 = pi044 & n5503;
  assign n7148 = ~n7146 & ~n7147;
  assign n7149 = n1521 & ~n7148;
  assign n7150 = ~n632 & ~n5228;
  assign n7151 = ~pi039 & ~n7150;
  assign n7152 = ~n793 & ~n5379;
  assign n7153 = pi039 & ~n7152;
  assign n7154 = ~n528 & ~n2329;
  assign n7155 = ~n7151 & n7154;
  assign n7156 = ~n7153 & n7155;
  assign n7157 = n6433 & ~n7156;
  assign n7158 = n1965 & n6332;
  assign n7159 = n492 & n6215;
  assign n7160 = ~n7158 & ~n7159;
  assign n7161 = pi065 & n1309;
  assign n7162 = ~n7160 & n7161;
  assign n7163 = ~n833 & ~n3008;
  assign n7164 = n6512 & ~n7163;
  assign n7165 = ~n1351 & ~n2291;
  assign n7166 = ~n2994 & n7165;
  assign n7167 = n7077 & ~n7166;
  assign n7168 = ~n7164 & ~n7167;
  assign n7169 = pi044 & ~n7168;
  assign n7170 = ~n2213 & ~n2898;
  assign n7171 = ~pi045 & ~n7170;
  assign n7172 = ~n2337 & n6447;
  assign n7173 = ~pi006 & n2685;
  assign n7174 = ~n2367 & ~n7173;
  assign n7175 = n2775 & n7174;
  assign n7176 = n6705 & n7175;
  assign n7177 = n5691 & n7176;
  assign n7178 = n7135 & ~n7177;
  assign n7179 = ~n1478 & n5663;
  assign n7180 = n329 & ~n7179;
  assign n7181 = n2779 & n2804;
  assign n7182 = ~pi029 & ~n7181;
  assign n7183 = pi039 & n3484;
  assign n7184 = n2392 & ~n3348;
  assign n7185 = n788 & ~n7184;
  assign n7186 = ~n2294 & n2932;
  assign n7187 = ~n5580 & ~n7186;
  assign n7188 = n1029 & ~n2723;
  assign n7189 = pi036 & n567;
  assign n7190 = ~n1317 & n7189;
  assign n7191 = n1298 & n7190;
  assign n7192 = ~n378 & ~n1971;
  assign n7193 = ~n2396 & ~n3175;
  assign n7194 = n5632 & ~n7183;
  assign n7195 = n7193 & n7194;
  assign n7196 = ~n4239 & n7192;
  assign n7197 = ~n6495 & n7187;
  assign n7198 = n7196 & n7197;
  assign n7199 = ~n2243 & n7195;
  assign n7200 = ~n2974 & ~n7185;
  assign n7201 = n7199 & n7200;
  assign n7202 = ~n2660 & n7198;
  assign n7203 = ~n2785 & n5667;
  assign n7204 = ~n6204 & ~n7191;
  assign n7205 = n7203 & n7204;
  assign n7206 = n7201 & n7202;
  assign n7207 = ~n3077 & n6035;
  assign n7208 = n7206 & n7207;
  assign n7209 = n2372 & n7205;
  assign n7210 = ~n3728 & ~n3826;
  assign n7211 = n5522 & n7066;
  assign n7212 = ~n7188 & n7211;
  assign n7213 = n7209 & n7210;
  assign n7214 = ~n2236 & n7208;
  assign n7215 = n2657 & ~n2844;
  assign n7216 = n7214 & n7215;
  assign n7217 = n7212 & n7213;
  assign n7218 = ~n7182 & n7217;
  assign n7219 = n3065 & n7216;
  assign n7220 = n5518 & n7219;
  assign n7221 = n7128 & n7218;
  assign n7222 = ~n7180 & n7221;
  assign n7223 = n7220 & n7222;
  assign n7224 = n6332 & ~n7223;
  assign n7225 = n771 & n1172;
  assign n7226 = ~n5367 & ~n7225;
  assign n7227 = n2282 & n7226;
  assign n7228 = n6504 & n7227;
  assign n7229 = ~n2829 & n7228;
  assign n7230 = n6660 & n7229;
  assign n7231 = n2381 & ~n7230;
  assign n7232 = ~n3068 & ~n5668;
  assign n7233 = n5577 & n7232;
  assign n7234 = n2942 & n7233;
  assign n7235 = n5563 & n7234;
  assign n7236 = n5557 & n7235;
  assign n7237 = n4405 & ~n7236;
  assign n7238 = ~n1440 & ~n1468;
  assign n7239 = ~n3637 & n7238;
  assign n7240 = n6431 & n7239;
  assign n7241 = n6380 & n7240;
  assign n7242 = n6305 & ~n7241;
  assign n7243 = n329 & n2381;
  assign n7244 = ~n3019 & n7243;
  assign n7245 = n2877 & ~n7244;
  assign n7246 = ~n7242 & n7245;
  assign n7247 = ~n7231 & n7246;
  assign n7248 = ~n7237 & n7247;
  assign n7249 = n5014 & ~n7248;
  assign n7250 = ~n7141 & ~n7172;
  assign n7251 = ~n7137 & n7250;
  assign n7252 = ~n7162 & n7251;
  assign n7253 = ~n7145 & ~n7149;
  assign n7254 = ~n7157 & n7253;
  assign n7255 = n7252 & n7254;
  assign n7256 = ~n7171 & n7255;
  assign n7257 = ~n7169 & n7256;
  assign n7258 = ~n7134 & n7257;
  assign n7259 = ~n7178 & n7258;
  assign n7260 = ~n7249 & n7259;
  assign po094 = n7224 | ~n7260;
  assign n7262 = n537 & n2035;
  assign n7263 = n1503 & ~n7262;
  assign n7264 = n1349 & n7263;
  assign n7265 = n3293 & n7264;
  assign po095 = ~n1320 | ~n7265;
  assign n7267 = n2893 & n3028;
  assign n7268 = n791 & ~n7267;
  assign n7269 = ~n2035 & ~n7161;
  assign n7270 = n2677 & ~n7269;
  assign n7271 = n1336 & n1473;
  assign n7272 = n1333 & n1376;
  assign n7273 = ~n2917 & ~n7270;
  assign n7274 = ~n7272 & n7273;
  assign n7275 = ~n7271 & n7274;
  assign n7276 = n7027 & n7275;
  assign po096 = n7268 | ~n7276;
  assign n7278 = n417 & n2999;
  assign n7279 = ~pi020 & ~n329;
  assign n7280 = n933 & ~n7279;
  assign n7281 = ~n2808 & ~n7280;
  assign n7282 = n1579 & ~n7281;
  assign n7283 = ~n7278 & ~n7282;
  assign n7284 = n2822 & n7283;
  assign n7285 = pi071 & ~n7284;
  assign n7286 = ~pi013 & n3798;
  assign n7287 = ~n2913 & ~n7286;
  assign n7288 = n1525 & n1955;
  assign n7289 = pi063 & n3212;
  assign n7290 = ~n5260 & ~n7288;
  assign n7291 = ~n6271 & ~n7289;
  assign n7292 = n7290 & n7291;
  assign n7293 = n2899 & n7292;
  assign n7294 = n7112 & n7293;
  assign n7295 = n7287 & n7294;
  assign po097 = n7285 | ~n7295;
  assign n7297 = ~n1464 & ~n1583;
  assign n7298 = n492 & ~n7297;
  assign n7299 = n329 & n906;
  assign n7300 = pi070 & ~n7284;
  assign n7301 = pi062 & n3212;
  assign n7302 = ~n6271 & ~n7301;
  assign n7303 = ~n7298 & n7302;
  assign n7304 = ~n2897 & n7303;
  assign n7305 = ~n7299 & n7304;
  assign po098 = n7300 | ~n7305;
  assign n7307 = pi061 & ~pi062;
  assign n7308 = n1168 & n7307;
  assign n7309 = n483 & n931;
  assign n7310 = ~n2671 & ~n7309;
  assign n7311 = n7308 & ~n7310;
  assign n7312 = n345 & n2656;
  assign n7313 = pi061 & n3212;
  assign n7314 = pi065 & ~n7284;
  assign n7315 = ~pi031 & pi062;
  assign n7316 = ~n2671 & ~n6273;
  assign n7317 = n7315 & ~n7316;
  assign n7318 = pi039 & n2411;
  assign n7319 = n1243 & n7318;
  assign n7320 = n938 & n7319;
  assign n7321 = n7315 & n7320;
  assign n7322 = n416 & n7308;
  assign n7323 = n7319 & n7322;
  assign n7324 = ~n7321 & ~n7323;
  assign n7325 = ~n7312 & ~n7313;
  assign n7326 = ~n2898 & n7325;
  assign n7327 = ~n2904 & n7326;
  assign n7328 = ~n7030 & n7327;
  assign n7329 = ~n7317 & n7324;
  assign n7330 = n7328 & n7329;
  assign n7331 = n7287 & ~n7311;
  assign n7332 = n7330 & n7331;
  assign po099 = n7314 | ~n7332;
  assign n7334 = pi049 & ~pi052;
  assign n7335 = n3602 & n7334;
  assign n7336 = pi015 & n4010;
  assign n7337 = ~n7335 & ~n7336;
  assign n7338 = n1596 & n3203;
  assign n7339 = ~pi106 & n4379;
  assign n7340 = n533 & ~n4537;
  assign n7341 = ~pi083 & n1228;
  assign n7342 = ~pi086 & n1965;
  assign n7343 = ~pi085 & n1030;
  assign n7344 = ~pi087 & n1306;
  assign n7345 = ~pi084 & n1338;
  assign n7346 = ~pi082 & n798;
  assign n7347 = ~pi081 & n330;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = pi045 & ~n7348;
  assign n7350 = ~n7341 & ~n7343;
  assign n7351 = ~n7345 & n7350;
  assign n7352 = ~n7342 & ~n7344;
  assign n7353 = n7351 & n7352;
  assign n7354 = ~n7349 & n7353;
  assign n7355 = n1836 & ~n7354;
  assign n7356 = pi029 & pi081;
  assign n7357 = ~pi029 & pi080;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = n2680 & n7358;
  assign n7360 = n2071 & n7359;
  assign n7361 = pi050 & ~pi051;
  assign n7362 = n4148 & n7361;
  assign n7363 = pi089 & ~n3795;
  assign n7364 = pi088 & n527;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = ~pi051 & ~n7365;
  assign n7367 = n875 & n3011;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = ~n7362 & n7368;
  assign n7370 = ~pi051 & ~pi077;
  assign n7371 = pi048 & n442;
  assign n7372 = n340 & n7371;
  assign po106 = n7370 & n7372;
  assign po102 = ~n7369 | po106;
  assign n7375 = n338 & n500;
  assign n7376 = ~pi062 & n7375;
  assign n7377 = ~n1595 & ~n6196;
  assign n7378 = ~n7340 & ~n7376;
  assign n7379 = n7377 & n7378;
  assign n7380 = ~n7338 & ~n7339;
  assign n7381 = n7379 & n7380;
  assign n7382 = ~n7360 & n7381;
  assign n7383 = n3263 & n7382;
  assign n7384 = ~n7355 & n7383;
  assign n7385 = n3694 & n7337;
  assign n7386 = n7384 & n7385;
  assign po101 = po102 | ~n7386;
  assign n7388 = pi015 & po106;
  assign n7389 = ~pi051 & n7363;
  assign n7390 = ~pi015 & n7362;
  assign n7391 = ~n876 & ~n7390;
  assign n7392 = ~n7388 & n7391;
  assign po103 = n7389 | ~n7392;
  assign n7394 = n442 & n7361;
  assign n7395 = n723 & n7394;
  assign po104 = n7366 | n7395;
  assign po105 = ~n7337 | ~n7369;
  assign n7398 = pi015 & n7362;
  assign n7399 = ~po106 & ~n7398;
  assign n7400 = n7337 & n7399;
  assign po107 = ~n7368 | ~n7400;
  assign n7402 = ~n2765 & ~n5162;
  assign po108 = ~n2852 | ~n7402;
  assign n7404 = n1699 & n4124;
  assign n7405 = ~n1749 & n4853;
  assign n7406 = n898 & ~n7405;
  assign n7407 = ~n1706 & ~n1719;
  assign n7408 = ~n2544 & ~n7404;
  assign n7409 = n7407 & n7408;
  assign n7410 = ~n7406 & n7409;
  assign n7411 = ~n2525 & n7410;
  assign n7412 = ~n4059 & ~n4796;
  assign n7413 = n1718 & ~n7412;
  assign n7414 = n1702 & n1990;
  assign n7415 = ~n1671 & ~n1700;
  assign n7416 = n3473 & ~n7415;
  assign n7417 = n330 & ~n3303;
  assign n7418 = n2604 & ~n7414;
  assign n7419 = ~n7413 & ~n7416;
  assign n7420 = ~n7417 & n7419;
  assign n7421 = n7418 & n7420;
  assign n7422 = n7411 & n7421;
  assign po114 = ~n6492 | ~n7422;
  assign n7424 = n2547 & ~n4556;
  assign n7425 = ~n4728 & n7424;
  assign n7426 = n2502 & n7425;
  assign po116 = n2574 | ~n7426;
  assign n7428 = ~pi029 & n1158;
  assign n7429 = n408 & ~n7428;
  assign n7430 = ~n750 & n7429;
  assign n7431 = ~n1766 & ~n3464;
  assign n7432 = ~po123 & ~n7430;
  assign po117 = ~n7431 | ~n7432;
  assign n7434 = ~n2038 & ~n2589;
  assign n7435 = n5952 & n7434;
  assign po118 = ~n2501 | ~n7435;
  assign n7437 = pi014 & ~n6864;
  assign n7438 = n1325 & n3295;
  assign po119 = n7437 | n7438;
  assign n7440 = ~n1719 & ~n2555;
  assign n7441 = n2526 & n6861;
  assign n7442 = n2605 & n7441;
  assign po120 = ~n7440 | ~n7442;
  assign po122 = n4047 | ~n7440;
  assign n7445 = n1234 & n1571;
  assign n7446 = ~n2094 & ~n7445;
  assign n7447 = ~pi019 & n414;
  assign n7448 = n1898 & ~n1999;
  assign n7449 = n7446 & n7448;
  assign n7450 = n3909 & n7449;
  assign n7451 = n6270 & ~n7447;
  assign n7452 = n7450 & n7451;
  assign po124 = n3739 | ~n7452;
  assign n7454 = n1702 & ~n1991;
  assign n7455 = ~pi023 & n4574;
  assign n7456 = ~pi015 & n2602;
  assign n7457 = n300 & n2051;
  assign n7458 = n381 & ~n391;
  assign n7459 = ~n394 & ~n7458;
  assign n7460 = n2301 & n4029;
  assign n7461 = ~pi122 & n404;
  assign n7462 = n345 & n550;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = n377 & ~n7463;
  assign n7465 = ~n7460 & ~n7464;
  assign n7466 = ~n4231 & n7465;
  assign n7467 = ~n7457 & n7466;
  assign n7468 = ~n6947 & ~n7455;
  assign n7469 = ~n7459 & n7468;
  assign n7470 = ~n3683 & n7467;
  assign n7471 = ~n7454 & ~n7456;
  assign n7472 = n7470 & n7471;
  assign n7473 = ~n383 & n7469;
  assign n7474 = n2500 & n7424;
  assign n7475 = n7473 & n7474;
  assign n7476 = n7410 & n7472;
  assign n7477 = n7475 & n7476;
  assign n7478 = n7452 & n7477;
  assign po125 = ~n2593 | ~n7478;
  assign n7480 = n653 & n4473;
  assign n7481 = ~n711 & ~n7480;
  assign n7482 = pi013 & ~n7481;
  assign n7483 = ~n3739 & ~n3906;
  assign n7484 = n1232 & n7483;
  assign n7485 = n5005 & n7484;
  assign po126 = n7482 | ~n7485;
  assign n7487 = ~pi023 & n2096;
  assign n7488 = pi065 & n1294;
  assign n7489 = n2567 & ~n7488;
  assign n7490 = n537 & ~n7489;
  assign n7491 = n798 & n2720;
  assign n7492 = n395 & n3537;
  assign n7493 = n585 & ~n1777;
  assign n7494 = n1833 & ~n7493;
  assign n7495 = n492 & ~n7494;
  assign n7496 = ~po072 & n7431;
  assign n7497 = ~n7487 & ~n7491;
  assign n7498 = n7496 & n7497;
  assign n7499 = n7440 & n7498;
  assign n7500 = ~n7482 & n7499;
  assign n7501 = n6858 & ~n7490;
  assign n7502 = n7492 & n7501;
  assign n7503 = n7500 & n7502;
  assign n7504 = n2613 & ~n7495;
  assign po127 = ~n7503 | ~n7504;
  assign n7506 = pi065 & n2590;
  assign po128 = n557 | n7506;
  assign n7508 = ~pi097 & pi098;
  assign n7509 = n2814 & n7508;
  assign n7510 = ~pi045 & n498;
  assign n7511 = pi045 & n833;
  assign n7512 = ~n7510 & ~n7511;
  assign n7513 = n832 & ~n7512;
  assign po129 = n7509 | n7513;
  assign n7515 = ~n1158 & n2860;
  assign n7516 = ~n1169 & ~n7515;
  assign n7517 = n2816 & n7508;
  assign n7518 = ~n1596 & ~n5397;
  assign n7519 = n3203 & ~n7518;
  assign n7520 = ~n1138 & n1150;
  assign n7521 = pi108 & n308;
  assign n7522 = n3103 & n7521;
  assign n7523 = ~n999 & n7522;
  assign n7524 = pi097 & n2814;
  assign n7525 = pi039 & n2698;
  assign n7526 = n7307 & n7320;
  assign n7527 = ~n7525 & ~n7526;
  assign n7528 = ~pi031 & ~n7527;
  assign n7529 = n329 & n814;
  assign n7530 = ~pi034 & n7375;
  assign n7531 = ~pi033 & n7530;
  assign n7532 = pi045 & ~n498;
  assign n7533 = ~pi045 & ~n833;
  assign n7534 = n832 & ~n7532;
  assign n7535 = ~n7533 & n7534;
  assign n7536 = n829 & n7510;
  assign n7537 = ~n7531 & ~n7536;
  assign n7538 = ~n7535 & n7537;
  assign n7539 = ~n7519 & ~n7523;
  assign n7540 = n7538 & n7539;
  assign n7541 = ~n7520 & n7540;
  assign n7542 = n7516 & ~n7517;
  assign n7543 = n7541 & n7542;
  assign n7544 = ~n7311 & ~n7528;
  assign n7545 = n7543 & n7544;
  assign n7546 = ~n2186 & ~n7529;
  assign n7547 = n7545 & n7546;
  assign n7548 = n2184 & n7547;
  assign n7549 = n3830 & ~n7524;
  assign po130 = ~n7548 | ~n7549;
  assign n7551 = pi045 & n829;
  assign n7552 = ~n834 & n7551;
  assign n7553 = n3099 & ~n5246;
  assign n7554 = ~pi045 & ~n2372;
  assign n7555 = n751 & n7521;
  assign n7556 = ~n999 & n1054;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = n3103 & ~n7557;
  assign n7559 = ~n2752 & n7016;
  assign n7560 = ~n1272 & ~n4765;
  assign n7561 = n4731 & n7560;
  assign n7562 = n7559 & n7561;
  assign n7563 = pi065 & ~n7562;
  assign n7564 = ~n766 & n3103;
  assign n7565 = ~n842 & ~n7564;
  assign n7566 = pi108 & ~n7565;
  assign n7567 = ~pi031 & n2671;
  assign n7568 = pi122 & n7307;
  assign n7569 = ~pi062 & ~n7568;
  assign n7570 = n7567 & ~n7569;
  assign n7571 = ~pi034 & n1595;
  assign n7572 = ~n7525 & ~n7571;
  assign n7573 = pi031 & ~n7572;
  assign n7574 = ~n1596 & ~n7375;
  assign n7575 = pi034 & ~n7574;
  assign n7576 = ~pi039 & n5495;
  assign n7577 = ~n1913 & ~n7576;
  assign n7578 = n4066 & n7577;
  assign n7579 = n2646 & ~n7578;
  assign n7580 = n572 & n867;
  assign n7581 = n408 & ~n1919;
  assign n7582 = ~n2677 & ~n7581;
  assign n7583 = ~n1306 & n7582;
  assign n7584 = n7488 & ~n7583;
  assign n7585 = ~pi031 & pi034;
  assign n7586 = n1599 & n7585;
  assign n7587 = ~n3010 & n6892;
  assign n7588 = ~n7077 & ~n7587;
  assign n7589 = n329 & ~n5502;
  assign n7590 = ~n879 & ~n7589;
  assign n7591 = ~n7588 & ~n7590;
  assign n7592 = pi033 & n7530;
  assign n7593 = pi097 & ~n2817;
  assign n7594 = pi051 & n829;
  assign n7595 = n874 & n7594;
  assign n7596 = ~n1133 & ~n7595;
  assign n7597 = ~n7592 & n7596;
  assign n7598 = ~n1993 & n7597;
  assign n7599 = ~n3107 & n7598;
  assign n7600 = ~n4745 & n7599;
  assign n7601 = ~n7593 & n7600;
  assign n7602 = pi062 & n6273;
  assign n7603 = ~n7307 & n7320;
  assign n7604 = n345 & n7309;
  assign n7605 = n7307 & n7604;
  assign n7606 = pi039 & ~n2700;
  assign n7607 = ~pi032 & ~n7606;
  assign n7608 = ~n2701 & n7607;
  assign n7609 = ~n7602 & ~n7608;
  assign n7610 = ~n7603 & n7609;
  assign n7611 = ~n7605 & n7610;
  assign n7612 = ~pi031 & ~n7611;
  assign n7613 = ~n6493 & ~n6802;
  assign n7614 = ~pi039 & ~n7613;
  assign n7615 = ~n1207 & ~n7586;
  assign n7616 = ~n1182 & n7615;
  assign n7617 = ~n2017 & ~n7580;
  assign n7618 = n7616 & n7617;
  assign n7619 = ~n7535 & ~n7552;
  assign n7620 = ~n7584 & n7619;
  assign n7621 = ~n2811 & n7618;
  assign n7622 = ~n7570 & ~n7575;
  assign n7623 = n7621 & n7622;
  assign n7624 = ~n1334 & n7620;
  assign n7625 = ~n7553 & ~n7573;
  assign n7626 = n7624 & n7625;
  assign n7627 = ~n846 & n7623;
  assign n7628 = ~n2185 & ~n7558;
  assign n7629 = n7627 & n7628;
  assign n7630 = ~n7554 & n7626;
  assign n7631 = ~n7563 & n7630;
  assign n7632 = n1454 & n7629;
  assign n7633 = ~n4223 & ~n7490;
  assign n7634 = ~n7566 & ~n7579;
  assign n7635 = n7633 & n7634;
  assign n7636 = n7631 & n7632;
  assign n7637 = ~n1737 & n2617;
  assign n7638 = ~n7015 & n7022;
  assign n7639 = ~n7591 & ~n7612;
  assign n7640 = n7638 & n7639;
  assign n7641 = n7636 & n7637;
  assign n7642 = ~n7614 & n7635;
  assign n7643 = n7641 & n7642;
  assign n7644 = n7640 & n7643;
  assign po131 = ~n7601 | ~n7644;
  assign n7646 = ~pi045 & ~n2378;
  assign n7647 = ~n802 & ~n1030;
  assign n7648 = ~n1305 & n7647;
  assign n7649 = n1301 & ~n7648;
  assign n7650 = ~n6188 & ~n7649;
  assign n7651 = ~n360 & ~n7650;
  assign n7652 = ~n330 & ~n1338;
  assign n7653 = ~n1964 & n7652;
  assign n7654 = n1301 & ~n7653;
  assign n7655 = ~n3818 & ~n5874;
  assign n7656 = pi067 & ~n7655;
  assign n7657 = ~pi066 & ~n783;
  assign n7658 = n328 & n7657;
  assign n7659 = n751 & n1054;
  assign n7660 = ~n344 & n2035;
  assign n7661 = n307 & n867;
  assign n7662 = ~pi058 & ~pi059;
  assign n7663 = n1623 & ~n7662;
  assign n7664 = ~n325 & ~n7663;
  assign n7665 = n329 & ~n7664;
  assign n7666 = ~n998 & ~n7659;
  assign n7667 = ~n5537 & ~n7660;
  assign n7668 = ~n7661 & n7667;
  assign n7669 = n7666 & n7668;
  assign n7670 = ~n7665 & n7669;
  assign n7671 = n3103 & ~n7670;
  assign n7672 = ~n3055 & ~n4169;
  assign n7673 = n537 & ~n7672;
  assign n7674 = n741 & n3103;
  assign n7675 = ~n869 & ~n7674;
  assign n7676 = pi108 & ~n7675;
  assign n7677 = pi104 & n2927;
  assign n7678 = ~pi061 & ~pi062;
  assign n7679 = n1168 & n7678;
  assign n7680 = n7309 & n7679;
  assign n7681 = ~pi088 & n527;
  assign n7682 = ~n880 & ~n3007;
  assign n7683 = ~pi039 & ~n7682;
  assign n7684 = n345 & n1268;
  assign n7685 = ~n3999 & ~n4765;
  assign n7686 = ~n7684 & n7685;
  assign n7687 = ~n1887 & n7686;
  assign n7688 = ~n4748 & n7687;
  assign n7689 = pi061 & ~n7688;
  assign n7690 = pi051 & ~n7365;
  assign n7691 = ~n7568 & ~n7678;
  assign n7692 = n7567 & ~n7691;
  assign n7693 = n4148 & ~n7361;
  assign n7694 = ~n329 & ~n1517;
  assign n7695 = n1915 & ~n7694;
  assign n7696 = ~pi048 & n442;
  assign n7697 = n340 & n7696;
  assign n7698 = ~n7106 & n7525;
  assign n7699 = ~pi045 & n2360;
  assign n7700 = n1145 & ~n1158;
  assign n7701 = n535 & n1837;
  assign n7702 = n345 & n1178;
  assign n7703 = n1270 & n7702;
  assign n7704 = ~pi039 & n3012;
  assign n7705 = pi039 & n1351;
  assign n7706 = n2036 & n2662;
  assign n7707 = pi122 & n1883;
  assign n7708 = pi034 & n1595;
  assign n7709 = pi074 & n432;
  assign n7710 = ~pi106 & n2703;
  assign n7711 = n1569 & n1571;
  assign n7712 = pi105 & n1445;
  assign n7713 = ~n1158 & n1175;
  assign n7714 = n829 & n833;
  assign n7715 = ~n7370 & n7372;
  assign n7716 = ~n1305 & ~n1308;
  assign n7717 = n1310 & ~n7716;
  assign n7718 = n7107 & ~n7606;
  assign n7719 = pi054 & n855;
  assign n7720 = ~n498 & ~n875;
  assign n7721 = n832 & ~n7720;
  assign n7722 = ~n3103 & ~n7429;
  assign n7723 = ~pi108 & ~n750;
  assign n7724 = ~n7722 & n7723;
  assign n7725 = ~pi040 & ~pi041;
  assign n7726 = n329 & n577;
  assign n7727 = ~n429 & ~n7726;
  assign n7728 = n1624 & ~n7725;
  assign n7729 = ~n7727 & n7728;
  assign n7730 = ~n740 & ~n1375;
  assign n7731 = n2880 & ~n7730;
  assign n7732 = ~n2674 & n5246;
  assign n7733 = n3869 & ~n7732;
  assign n7734 = pi039 & n4631;
  assign n7735 = ~pi031 & ~pi062;
  assign n7736 = n7604 & n7735;
  assign n7737 = ~n329 & ~n1965;
  assign n7738 = ~n344 & ~n7737;
  assign n7739 = ~n537 & ~n7738;
  assign n7740 = n1294 & ~n7739;
  assign n7741 = pi006 & n2684;
  assign n7742 = ~n5690 & ~n7741;
  assign n7743 = ~pi122 & n798;
  assign n7744 = ~n7742 & n7743;
  assign n7745 = ~n2756 & ~n7744;
  assign n7746 = ~n7740 & n7745;
  assign n7747 = pi061 & ~n7746;
  assign n7748 = ~n474 & n6671;
  assign n7749 = n1523 & ~n7727;
  assign n7750 = ~n3338 & ~n7749;
  assign n7751 = ~n7662 & ~n7750;
  assign n7752 = n763 & n3103;
  assign n7753 = ~n3324 & ~n7752;
  assign n7754 = ~pi124 & ~n7753;
  assign n7755 = n1599 & n3203;
  assign n7756 = pi031 & n7320;
  assign n7757 = ~n1334 & ~n7038;
  assign n7758 = ~n865 & ~n7681;
  assign n7759 = ~n7711 & ~n7755;
  assign n7760 = n7758 & n7759;
  assign n7761 = ~n7262 & ~n7693;
  assign n7762 = ~n7697 & ~n7703;
  assign n7763 = ~n7704 & ~n7705;
  assign n7764 = ~n7707 & ~n7712;
  assign n7765 = ~n7713 & ~n7714;
  assign n7766 = n7764 & n7765;
  assign n7767 = n7762 & n7763;
  assign n7768 = n7760 & n7761;
  assign n7769 = ~n2813 & ~n3843;
  assign n7770 = ~n7695 & ~n7706;
  assign n7771 = ~n7708 & ~n7710;
  assign n7772 = ~n7715 & ~n7717;
  assign n7773 = n7771 & n7772;
  assign n7774 = n7769 & n7770;
  assign n7775 = n7767 & n7768;
  assign n7776 = ~n1195 & n7766;
  assign n7777 = ~n1889 & ~n2382;
  assign n7778 = ~n2665 & ~n3696;
  assign n7779 = ~n4752 & ~n7692;
  assign n7780 = ~n7698 & ~n7709;
  assign n7781 = ~n7721 & ~n7733;
  assign n7782 = n7780 & n7781;
  assign n7783 = n7778 & n7779;
  assign n7784 = n7776 & n7777;
  assign n7785 = n7774 & n7775;
  assign n7786 = ~n2659 & n7773;
  assign n7787 = ~n5331 & ~n7335;
  assign n7788 = ~n7699 & ~n7700;
  assign n7789 = ~n7701 & ~n7718;
  assign n7790 = ~n7719 & ~n7724;
  assign n7791 = ~n7729 & ~n7731;
  assign n7792 = ~n7756 & n7791;
  assign n7793 = n7789 & n7790;
  assign n7794 = n7787 & n7788;
  assign n7795 = n7785 & n7786;
  assign n7796 = n7783 & n7784;
  assign n7797 = ~n2503 & n7782;
  assign n7798 = ~n2883 & ~n3793;
  assign n7799 = n7324 & ~n7676;
  assign n7800 = ~n7677 & ~n7680;
  assign n7801 = ~n7748 & ~n7754;
  assign n7802 = n7757 & n7801;
  assign n7803 = n7799 & n7800;
  assign n7804 = n7797 & n7798;
  assign n7805 = n7795 & n7796;
  assign n7806 = n7793 & n7794;
  assign n7807 = n850 & n7792;
  assign n7808 = n4985 & ~n7646;
  assign n7809 = ~n7654 & ~n7656;
  assign n7810 = ~n7671 & ~n7673;
  assign n7811 = ~n7736 & ~n7747;
  assign n7812 = ~n7751 & n7811;
  assign n7813 = n7809 & n7810;
  assign n7814 = n7807 & n7808;
  assign n7815 = n7805 & n7806;
  assign n7816 = n7803 & n7804;
  assign n7817 = n4071 & n7802;
  assign n7818 = ~n7658 & ~n7689;
  assign n7819 = ~n7690 & ~n7734;
  assign n7820 = n7818 & n7819;
  assign n7821 = n7816 & n7817;
  assign n7822 = n7814 & n7815;
  assign n7823 = n7812 & n7813;
  assign n7824 = ~n1882 & n2187;
  assign n7825 = n5775 & ~n7651;
  assign n7826 = n7824 & n7825;
  assign n7827 = n7822 & n7823;
  assign n7828 = n7820 & n7821;
  assign n7829 = n7827 & n7828;
  assign n7830 = ~n7683 & n7826;
  assign n7831 = n7829 & n7830;
  assign po132 = ~n7601 | ~n7831;
  assign n7833 = ~n2367 & ~n2920;
  assign n7834 = n2795 & n7833;
  assign n7835 = n5041 & n7834;
  assign n7836 = n329 & ~n7835;
  assign n7837 = ~pi015 & n2063;
  assign n7838 = n450 & n960;
  assign n7839 = n609 & n693;
  assign n7840 = ~n1702 & ~n3852;
  assign n7841 = n620 & ~n7840;
  assign n7842 = ~n7838 & ~n7841;
  assign n7843 = ~n7839 & n7842;
  assign n7844 = n290 & ~n7843;
  assign n7845 = n346 & n599;
  assign n7846 = ~n4214 & ~n7845;
  assign n7847 = n410 & ~n7846;
  assign n7848 = ~n5879 & ~n6272;
  assign n7849 = pi018 & ~n7848;
  assign n7850 = n593 & ~n4469;
  assign n7851 = n386 & n1380;
  assign n7852 = ~pi022 & n931;
  assign n7853 = ~n1388 & ~n7851;
  assign n7854 = ~n7852 & n7853;
  assign n7855 = n293 & ~n7854;
  assign n7856 = ~n3484 & ~n7186;
  assign n7857 = ~n3058 & n7856;
  assign n7858 = ~n3062 & n7857;
  assign n7859 = ~n7850 & n7858;
  assign n7860 = ~n7855 & n7859;
  assign n7861 = ~n474 & ~n7860;
  assign n7862 = n415 & ~n2039;
  assign n7863 = n2588 & n7862;
  assign n7864 = ~n467 & ~n683;
  assign n7865 = n302 & ~n7864;
  assign n7866 = ~pi015 & n1744;
  assign n7867 = ~n665 & ~n863;
  assign n7868 = ~n7866 & n7867;
  assign n7869 = n442 & ~n7868;
  assign n7870 = ~n7865 & ~n7869;
  assign n7871 = ~pi011 & ~n7870;
  assign n7872 = n2989 & n4036;
  assign n7873 = n345 & ~n7872;
  assign n7874 = ~pi105 & n1445;
  assign n7875 = ~n381 & n406;
  assign n7876 = n1917 & ~n7875;
  assign n7877 = n492 & ~n7876;
  assign n7878 = ~n2001 & ~n2335;
  assign n7879 = n335 & ~n7878;
  assign n7880 = n3011 & n7510;
  assign n7881 = ~n750 & n1093;
  assign n7882 = n756 & ~n1398;
  assign n7883 = ~n479 & ~n549;
  assign n7884 = n2075 & n7883;
  assign n7885 = n4427 & n7576;
  assign n7886 = ~n3590 & ~n3624;
  assign n7887 = ~pi018 & ~n7886;
  assign n7888 = ~n1095 & ~n1337;
  assign n7889 = n1336 & ~n7888;
  assign n7890 = n962 & n3473;
  assign n7891 = n1517 & n1521;
  assign n7892 = ~n368 & ~n4124;
  assign n7893 = n3295 & ~n7892;
  assign n7894 = n486 & n1688;
  assign n7895 = n1066 & n1076;
  assign n7896 = pi015 & n1760;
  assign n7897 = ~n485 & n1873;
  assign n7898 = ~n5885 & ~n7897;
  assign n7899 = n1081 & ~n7898;
  assign n7900 = pi023 & n1363;
  assign n7901 = n1362 & ~n7900;
  assign n7902 = n1590 & ~n7901;
  assign n7903 = n389 & n1047;
  assign n7904 = pi019 & n7903;
  assign n7905 = ~n405 & ~n1397;
  assign n7906 = n453 & ~n7905;
  assign n7907 = n375 & n416;
  assign n7908 = ~n2001 & ~n7907;
  assign n7909 = ~n7906 & n7908;
  assign n7910 = n529 & ~n7909;
  assign n7911 = ~n368 & ~n589;
  assign n7912 = n966 & ~n7911;
  assign n7913 = ~n3893 & ~n7912;
  assign n7914 = ~pi006 & ~n7913;
  assign n7915 = ~n644 & ~n1387;
  assign n7916 = n1047 & ~n7915;
  assign n7917 = ~n1016 & ~n1090;
  assign n7918 = pi006 & ~n7917;
  assign n7919 = pi029 & ~n879;
  assign n7920 = n7077 & ~n7919;
  assign n7921 = ~n7590 & n7920;
  assign n7922 = ~n6493 & ~n6803;
  assign n7923 = ~pi039 & ~n7922;
  assign n7924 = ~n360 & n6675;
  assign n7925 = n2945 & n2947;
  assign n7926 = n883 & n1243;
  assign n7927 = ~n6149 & ~n7926;
  assign n7928 = ~n3084 & n7927;
  assign n7929 = n361 & ~n7928;
  assign n7930 = ~n7924 & ~n7925;
  assign n7931 = ~n7929 & n7930;
  assign n7932 = ~n1166 & ~n2504;
  assign n7933 = ~n2333 & ~n7882;
  assign n7934 = ~n7884 & n7933;
  assign n7935 = ~n341 & n7932;
  assign n7936 = ~n4576 & ~n7874;
  assign n7937 = ~n7879 & ~n7880;
  assign n7938 = ~n7894 & ~n7904;
  assign n7939 = n7937 & n7938;
  assign n7940 = n7935 & n7936;
  assign n7941 = ~n1642 & n7934;
  assign n7942 = ~n1719 & ~n1856;
  assign n7943 = ~n3000 & ~n3695;
  assign n7944 = ~n7881 & ~n7885;
  assign n7945 = ~n7899 & ~n7910;
  assign n7946 = n7944 & n7945;
  assign n7947 = n7942 & n7943;
  assign n7948 = n7940 & n7941;
  assign n7949 = ~n612 & n7939;
  assign n7950 = n2315 & ~n2404;
  assign n7951 = ~n2898 & ~n3454;
  assign n7952 = ~n3480 & ~n6890;
  assign n7953 = ~n7459 & ~n7837;
  assign n7954 = ~n7893 & ~n7895;
  assign n7955 = ~n7896 & ~n7902;
  assign n7956 = ~n7914 & ~n7918;
  assign n7957 = n7955 & n7956;
  assign n7958 = n7953 & n7954;
  assign n7959 = n7951 & n7952;
  assign n7960 = n7949 & n7950;
  assign n7961 = n7947 & n7948;
  assign n7962 = ~n441 & n7946;
  assign n7963 = n712 & n1374;
  assign n7964 = ~n2927 & n2959;
  assign n7965 = n4643 & ~n4983;
  assign n7966 = n5324 & ~n7847;
  assign n7967 = ~n7849 & ~n7877;
  assign n7968 = ~n7890 & ~n7891;
  assign n7969 = ~n7916 & n7968;
  assign n7970 = n7966 & n7967;
  assign n7971 = n7964 & n7965;
  assign n7972 = n7962 & n7963;
  assign n7973 = n7960 & n7961;
  assign n7974 = n7958 & n7959;
  assign n7975 = n1734 & n7957;
  assign n7976 = n2749 & n3616;
  assign n7977 = n4836 & n7757;
  assign n7978 = ~n7844 & n7977;
  assign n7979 = n7975 & n7976;
  assign n7980 = n7973 & n7974;
  assign n7981 = n7971 & n7972;
  assign n7982 = n7969 & n7970;
  assign n7983 = n2766 & n3575;
  assign n7984 = n3987 & n4052;
  assign n7985 = n4432 & ~n4917;
  assign n7986 = n5037 & n5170;
  assign n7987 = ~n5425 & ~n5781;
  assign n7988 = ~n6766 & ~n7873;
  assign n7989 = ~n7887 & ~n7889;
  assign n7990 = n7931 & n7989;
  assign n7991 = n7987 & n7988;
  assign n7992 = n7985 & n7986;
  assign n7993 = n7983 & n7984;
  assign n7994 = n7981 & n7982;
  assign n7995 = n7979 & n7980;
  assign n7996 = n1509 & n7978;
  assign n7997 = n1575 & n3535;
  assign n7998 = n5265 & ~n7871;
  assign n7999 = n7997 & n7998;
  assign n8000 = n7995 & n7996;
  assign n8001 = n7993 & n7994;
  assign n8002 = n7991 & n7992;
  assign n8003 = n3291 & n7990;
  assign n8004 = n4187 & n5269;
  assign n8005 = ~n7861 & ~n7921;
  assign n8006 = n8004 & n8005;
  assign n8007 = n8002 & n8003;
  assign n8008 = n8000 & n8001;
  assign n8009 = n1312 & n7999;
  assign n8010 = n3323 & n5992;
  assign n8011 = n8009 & n8010;
  assign n8012 = n8007 & n8008;
  assign n8013 = n2742 & n8006;
  assign n8014 = n2984 & ~n3014;
  assign n8015 = n4235 & n4764;
  assign n8016 = n4928 & n5759;
  assign n8017 = ~n7923 & n8016;
  assign n8018 = n8014 & n8015;
  assign n8019 = n8012 & n8013;
  assign n8020 = n2872 & n8011;
  assign n8021 = ~n7836 & n7863;
  assign n8022 = n8020 & n8021;
  assign n8023 = n8018 & n8019;
  assign n8024 = n7020 & n8017;
  assign n8025 = n8023 & n8024;
  assign n8026 = n2823 & n8022;
  assign po133 = ~n8025 | ~n8026;
  assign n8028 = n1247 & n1375;
  assign n8029 = n2667 & ~n8028;
  assign n8030 = n2609 & n8029;
  assign n8031 = ~n2647 & n8030;
  assign po134 = n1222 | ~n8031;
  assign n8033 = ~pi122 & n2798;
  assign n8034 = n592 & n8033;
  assign n8035 = ~pi013 & n2034;
  assign n8036 = n515 & n4172;
  assign n8037 = n1375 & ~n3257;
  assign n8038 = n2539 & n8037;
  assign n8039 = ~n1222 & ~n1281;
  assign n8040 = n5254 & n8039;
  assign n8041 = n2726 & n8040;
  assign n8042 = ~n8034 & ~n8036;
  assign n8043 = ~n2670 & n8042;
  assign n8044 = ~n8038 & n8043;
  assign n8045 = ~n8035 & n8044;
  assign n8046 = n4991 & ~n7271;
  assign n8047 = n8045 & n8046;
  assign n8048 = n8041 & n8047;
  assign po138 = ~n8031 | ~n8048;
  assign n8050 = ~po002 & n4478;
  assign n8051 = n4920 & n8050;
  assign n8052 = ~n5585 & n8051;
  assign n8053 = ~n1328 & ~n2769;
  assign n8054 = n4766 & n8053;
  assign n8055 = n791 & ~n8054;
  assign n8056 = n2846 & n5330;
  assign n8057 = ~n937 & ~n1259;
  assign n8058 = ~n3081 & n8057;
  assign n8059 = n361 & ~n8058;
  assign n8060 = pi001 & n1397;
  assign n8061 = ~n5528 & ~n8060;
  assign n8062 = n1385 & ~n8061;
  assign n8063 = ~pi003 & ~n3463;
  assign n8064 = n2650 & n8041;
  assign n8065 = n8030 & n8064;
  assign n8066 = ~pi023 & n2389;
  assign n8067 = ~pi019 & n7903;
  assign n8068 = pi022 & n1591;
  assign n8069 = ~n2077 & ~n2411;
  assign n8070 = n1712 & ~n8069;
  assign n8071 = ~n584 & n1368;
  assign n8072 = ~n1416 & ~n8071;
  assign n8073 = n442 & ~n8072;
  assign n8074 = ~n883 & ~n1027;
  assign n8075 = n1380 & ~n8074;
  assign n8076 = ~n1384 & ~n8075;
  assign n8077 = ~n3493 & n8076;
  assign n8078 = pi023 & n1385;
  assign n8079 = ~n8077 & n8078;
  assign n8080 = n3483 & ~n8067;
  assign n8081 = ~n8068 & n8080;
  assign n8082 = ~n8070 & n8081;
  assign n8083 = n2403 & n8082;
  assign n8084 = n5400 & ~n8066;
  assign n8085 = n8083 & n8084;
  assign n8086 = ~n8073 & ~n8079;
  assign n8087 = n8085 & n8086;
  assign n8088 = ~n2799 & ~n8063;
  assign n8089 = ~n8056 & n8088;
  assign n8090 = ~n8062 & n8089;
  assign n8091 = ~n8059 & n8090;
  assign n8092 = ~n1474 & n4588;
  assign n8093 = ~n8055 & n8092;
  assign n8094 = n8087 & n8091;
  assign n8095 = n8093 & n8094;
  assign n8096 = n8052 & n8095;
  assign n8097 = n3755 & n8096;
  assign po139 = ~n8065 | ~n8097;
  assign n8099 = n928 & ~n2951;
  assign n8100 = n699 & n1975;
  assign n8101 = ~n3734 & ~n4239;
  assign n8102 = ~n8100 & n8101;
  assign n8103 = n7032 & n8102;
  assign n8104 = ~n2776 & n8103;
  assign n8105 = n4491 & n8104;
  assign n8106 = n8065 & n8105;
  assign n8107 = n2342 & ~n8099;
  assign n8108 = n7060 & n8107;
  assign n8109 = n8106 & n8108;
  assign n8110 = n1071 & n1275;
  assign n8111 = n2257 & ~n8110;
  assign n8112 = n3801 & n8111;
  assign n8113 = n293 & ~n8112;
  assign n8114 = ~pi003 & n3460;
  assign n8115 = n592 & n1868;
  assign n8116 = ~n2323 & ~n8114;
  assign n8117 = ~n8115 & n8116;
  assign n8118 = pi122 & ~n8117;
  assign n8119 = n6202 & n7187;
  assign n8120 = n2292 & n8119;
  assign n8121 = n6190 & ~n8118;
  assign n8122 = n8120 & n8121;
  assign n8123 = ~n8113 & n8122;
  assign n8124 = ~n360 & ~n8123;
  assign n8125 = n929 & n1243;
  assign n8126 = ~n364 & ~n8125;
  assign n8127 = ~n4267 & n8126;
  assign n8128 = ~pi018 & ~n8127;
  assign n8129 = ~n381 & ~n2876;
  assign n8130 = pi022 & n2785;
  assign n8131 = n376 & n8060;
  assign n8132 = ~n1506 & ~n8131;
  assign n8133 = ~n8130 & n8132;
  assign n8134 = ~pi122 & ~n8133;
  assign n8135 = n551 & ~n4000;
  assign n8136 = n725 & n2947;
  assign n8137 = n8072 & ~n8136;
  assign n8138 = pi012 & ~n8137;
  assign n8139 = n550 & n993;
  assign n8140 = n377 & n7461;
  assign n8141 = n1969 & n3494;
  assign n8142 = ~n8139 & ~n8140;
  assign n8143 = ~n2079 & n8142;
  assign n8144 = ~n2327 & n8143;
  assign n8145 = ~n3893 & ~n4270;
  assign n8146 = ~n8135 & n8145;
  assign n8147 = n8144 & n8146;
  assign n8148 = ~n2389 & ~n4579;
  assign n8149 = ~n8129 & ~n8141;
  assign n8150 = n8148 & n8149;
  assign n8151 = ~n1429 & n8147;
  assign n8152 = n8150 & n8151;
  assign n8153 = n1068 & n2960;
  assign n8154 = ~n4457 & ~n8128;
  assign n8155 = n8153 & n8154;
  assign n8156 = n2874 & n8152;
  assign n8157 = n4991 & ~n8134;
  assign n8158 = ~n8138 & n8157;
  assign n8159 = n8155 & n8156;
  assign n8160 = n8158 & n8159;
  assign n8161 = n8052 & ~n8124;
  assign n8162 = n8160 & n8161;
  assign n8163 = n2983 & n8162;
  assign po140 = ~n8109 | ~n8163;
  assign n8165 = n1064 & n1539;
  assign n8166 = n2259 & ~n8165;
  assign n8167 = n3092 & n8166;
  assign n8168 = n293 & ~n8167;
  assign n8169 = ~n3046 & ~n5633;
  assign n8170 = ~n1394 & n8169;
  assign n8171 = n2247 & n8170;
  assign n8172 = ~n8168 & n8171;
  assign n8173 = ~n360 & ~n8172;
  assign n8174 = n1969 & n2359;
  assign n8175 = n509 & n1590;
  assign n8176 = ~n2276 & ~n8175;
  assign n8177 = n361 & ~n8176;
  assign n8178 = n361 & n1049;
  assign n8179 = ~n7845 & ~n8178;
  assign n8180 = n417 & ~n8179;
  assign n8181 = ~n506 & ~n8178;
  assign n8182 = n933 & ~n8181;
  assign n8183 = n1368 & ~n2392;
  assign n8184 = ~pi020 & n8056;
  assign n8185 = pi022 & n641;
  assign n8186 = ~n792 & ~n8185;
  assign n8187 = ~n1519 & ~n2343;
  assign n8188 = n2092 & ~n8187;
  assign n8189 = n404 & n2296;
  assign n8190 = n306 & n2263;
  assign n8191 = n484 & n1366;
  assign n8192 = ~n6675 & ~n8189;
  assign n8193 = ~n8190 & n8192;
  assign n8194 = ~n8191 & n8193;
  assign n8195 = ~n474 & ~n8194;
  assign n8196 = ~pi004 & n2933;
  assign n8197 = ~n954 & ~n8196;
  assign n8198 = n453 & ~n8197;
  assign n8199 = ~n2303 & ~n4825;
  assign n8200 = ~n8198 & n8199;
  assign n8201 = ~n2389 & ~n2799;
  assign n8202 = n2949 & n4221;
  assign n8203 = ~n4999 & ~n8174;
  assign n8204 = ~n8183 & n8203;
  assign n8205 = n8201 & n8202;
  assign n8206 = ~n4593 & n8200;
  assign n8207 = ~n8180 & ~n8182;
  assign n8208 = ~n8184 & n8186;
  assign n8209 = ~n8188 & ~n8195;
  assign n8210 = n8208 & n8209;
  assign n8211 = n8206 & n8207;
  assign n8212 = n8204 & n8205;
  assign n8213 = ~n5424 & n8212;
  assign n8214 = n8210 & n8211;
  assign n8215 = n1430 & n8050;
  assign n8216 = ~n8177 & n8215;
  assign n8217 = n8213 & n8214;
  assign n8218 = n2968 & n8217;
  assign n8219 = n8216 & n8218;
  assign n8220 = n2984 & n8219;
  assign n8221 = n4216 & ~n8173;
  assign n8222 = n8220 & n8221;
  assign po141 = ~n8109 | ~n8222;
  assign n8224 = n1244 & n6894;
  assign n8225 = ~n2258 & n8058;
  assign n8226 = n8176 & n8225;
  assign n8227 = n361 & ~n8226;
  assign n8228 = ~n314 & ~n2066;
  assign n8229 = n954 & n8228;
  assign n8230 = pi014 & n4008;
  assign n8231 = n589 & n966;
  assign n8232 = n717 & n8178;
  assign n8233 = n1368 & ~n2390;
  assign n8234 = ~n444 & ~n725;
  assign n8235 = n314 & ~n8234;
  assign n8236 = ~n8233 & ~n8235;
  assign n8237 = n493 & ~n8236;
  assign n8238 = ~n360 & n717;
  assign n8239 = ~n1519 & ~n8238;
  assign n8240 = n2092 & ~n8239;
  assign n8241 = ~n993 & ~n4265;
  assign n8242 = n1397 & ~n8241;
  assign n8243 = n389 & n485;
  assign n8244 = n3247 & n8243;
  assign n8245 = ~n2774 & ~n3905;
  assign n8246 = ~n6180 & n8245;
  assign n8247 = n791 & ~n8246;
  assign n8248 = n1712 & n3628;
  assign n8249 = n906 & n1473;
  assign n8250 = n386 & n1969;
  assign n8251 = ~n8229 & ~n8231;
  assign n8252 = ~n8242 & ~n8244;
  assign n8253 = n8251 & n8252;
  assign n8254 = ~n4220 & ~n8230;
  assign n8255 = n8253 & n8254;
  assign n8256 = ~n8224 & ~n8232;
  assign n8257 = ~n8248 & ~n8250;
  assign n8258 = n8256 & n8257;
  assign n8259 = n8186 & n8255;
  assign n8260 = ~n8240 & n8259;
  assign n8261 = ~n8237 & n8258;
  assign n8262 = ~n8247 & n8261;
  assign n8263 = n3729 & n8260;
  assign n8264 = n7931 & n8263;
  assign n8265 = n1454 & n8262;
  assign n8266 = n4589 & n8051;
  assign n8267 = n8087 & ~n8227;
  assign n8268 = ~n8249 & n8267;
  assign n8269 = n8265 & n8266;
  assign n8270 = n3752 & n8264;
  assign n8271 = n8269 & n8270;
  assign po142 = ~n8268 | ~n8271;
  assign n8273 = ~n2244 & n2784;
  assign n8274 = ~pi122 & ~n8273;
  assign n8275 = n938 & ~n2271;
  assign n8276 = ~n1973 & ~n3726;
  assign n8277 = ~n7111 & ~n8034;
  assign n8278 = n8276 & n8277;
  assign n8279 = ~n2344 & n8278;
  assign n8280 = n796 & n2907;
  assign n8281 = ~n4477 & n8280;
  assign n8282 = ~n2305 & n8279;
  assign n8283 = n2673 & n2802;
  assign n8284 = ~n3728 & ~n7075;
  assign n8285 = n8283 & n8284;
  assign n8286 = n8281 & n8282;
  assign n8287 = ~n2991 & n3050;
  assign n8288 = ~n4161 & ~n8274;
  assign n8289 = ~n8275 & n8288;
  assign n8290 = n8286 & n8287;
  assign n8291 = n8285 & n8290;
  assign n8292 = n3318 & n8289;
  assign n8293 = n8291 & n8292;
  assign n8294 = n3098 & n8293;
  assign n8295 = n5264 & n8294;
  assign n8296 = n2987 & n8295;
  assign po143 = ~n8106 | ~n8296;
  assign n8298 = n1151 & ~n2854;
  assign n8299 = ~n1138 & ~n8298;
  assign n8300 = n2663 & n2758;
  assign n8301 = n2095 & n7033;
  assign n8302 = n791 & ~n2893;
  assign n8303 = n2743 & ~n3100;
  assign n8304 = ~n2017 & ~n7445;
  assign n8305 = n2676 & n8304;
  assign n8306 = ~n2710 & ~n8300;
  assign n8307 = n8305 & n8306;
  assign n8308 = n1209 & n8307;
  assign n8309 = n7516 & ~n8303;
  assign n8310 = n8308 & n8309;
  assign n8311 = n2750 & n2924;
  assign n8312 = n3108 & ~n8299;
  assign n8313 = n8301 & n8312;
  assign n8314 = n8310 & n8311;
  assign n8315 = n8313 & n8314;
  assign po144 = n8302 | ~n8315;
  assign n8317 = n1183 & ~n4448;
  assign n8318 = n1198 & n8317;
  assign n8319 = ~n1272 & ~n2993;
  assign n8320 = ~n2688 & n8319;
  assign n8321 = n2363 & n8320;
  assign n8322 = ~n4748 & n7559;
  assign n8323 = n8321 & n8322;
  assign po145 = ~n8318 | ~n8323;
  assign n8325 = n2684 & n2901;
  assign n8326 = n1440 & n4261;
  assign n8327 = ~n2756 & ~n8326;
  assign n8328 = ~n8325 & n8327;
  assign n8329 = ~n5268 & n8328;
  assign po146 = n2881 | ~n8329;
  assign n8331 = n1375 & ~n3027;
  assign n8332 = ~n5331 & ~n8331;
  assign po147 = po108 | ~n8332;
  assign n8334 = pi020 & n3901;
  assign n8335 = ~n1885 & ~n7404;
  assign n8336 = ~n775 & n6194;
  assign n8337 = n798 & ~n8336;
  assign n8338 = n601 & n604;
  assign n8339 = ~n2678 & ~n8338;
  assign n8340 = ~n8334 & n8339;
  assign n8341 = n8335 & n8340;
  assign n8342 = n4729 & ~n4811;
  assign n8343 = ~n8337 & n8342;
  assign n8344 = n8341 & n8343;
  assign po151 = n2574 | ~n8344;
  assign n8346 = n537 & n3055;
  assign n8347 = ~n6947 & ~n6954;
  assign n8348 = ~n8346 & n8347;
  assign po152 = po122 | ~n8348;
  assign n8350 = ~n2498 & ~n6162;
  assign n8351 = n1763 & ~n8350;
  assign n8352 = ~n2094 & ~n4556;
  assign n8353 = ~n8351 & n8352;
  assign n8354 = ~n711 & n8353;
  assign n8355 = ~n2495 & ~n3464;
  assign n8356 = n8354 & n8355;
  assign n8357 = ~n7454 & n8356;
  assign n8358 = n7411 & n8357;
  assign n8359 = n7492 & n8358;
  assign n8360 = n5154 & n8359;
  assign po153 = ~n2607 | ~n8360;
  assign n8362 = ~pi023 & ~n1423;
  assign n8363 = ~n1523 & ~n8362;
  assign n8364 = n6737 & ~n8363;
  assign n8365 = ~n337 & ~n370;
  assign n8366 = n744 & ~n8365;
  assign n8367 = ~n2396 & ~n8366;
  assign n8368 = ~n360 & ~n8367;
  assign n8369 = n2856 & ~n4417;
  assign n8370 = n5596 & ~n8369;
  assign n8371 = n2229 & n3267;
  assign n8372 = n596 & n1049;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n1261 & n8373;
  assign n8375 = n646 & n6892;
  assign n8376 = ~n8374 & n8375;
  assign n8377 = ~n1166 & ~n4409;
  assign n8378 = n2020 & n8377;
  assign n8379 = ~pi056 & ~n8378;
  assign n8380 = ~n1201 & ~n1221;
  assign n8381 = ~n5597 & ~n8380;
  assign n8382 = ~n775 & ~n6193;
  assign n8383 = n1228 & ~n8382;
  assign n8384 = n2365 & ~n2782;
  assign n8385 = ~n1281 & ~n6196;
  assign n8386 = ~n1995 & ~n2589;
  assign n8387 = n8385 & n8386;
  assign n8388 = ~n8364 & ~n8368;
  assign n8389 = n8387 & n8388;
  assign n8390 = ~n1456 & n5607;
  assign n8391 = n8389 & n8390;
  assign n8392 = n8318 & n8391;
  assign n8393 = ~n8376 & ~n8379;
  assign n8394 = ~n8381 & ~n8383;
  assign n8395 = n8393 & n8394;
  assign n8396 = ~n8370 & n8392;
  assign n8397 = n8395 & n8396;
  assign n8398 = ~n8384 & n8397;
  assign n8399 = n6930 & n8398;
  assign n8400 = n5947 & n8399;
  assign n8401 = ~n6701 & n8400;
  assign n8402 = ~n6883 & n8401;
  assign po154 = ~n6912 | ~n8402;
  assign n8404 = ~n1897 & n7446;
  assign n8405 = n2591 & n8404;
  assign n8406 = ~n4728 & n8405;
  assign n8407 = n8335 & n8406;
  assign po155 = ~n7863 | ~n8407;
  assign n8409 = n1233 & n8301;
  assign po156 = ~n2870 | ~n8409;
  assign n8411 = n991 & ~n1000;
  assign n8412 = ~n990 & ~n8411;
  assign n8413 = ~n5612 & ~n8412;
  assign n8414 = ~pi108 & ~n8413;
  assign n8415 = n3828 & ~n7919;
  assign n8416 = ~n376 & ~n1053;
  assign n8417 = n1020 & ~n8416;
  assign n8418 = n492 & n814;
  assign n8419 = ~n836 & ~n8417;
  assign n8420 = n877 & n8419;
  assign n8421 = ~n8414 & ~n8418;
  assign n8422 = n8420 & n8421;
  assign po158 = n8415 | ~n8422;
  assign n8424 = n330 & n7657;
  assign po159 = n1321 | n8424;
  assign po005 = 1'b0;
  assign po006 = 1'b0;
  assign po007 = 1'b0;
  assign po045 = 1'b0;
  assign po049 = 1'b0;
  assign po085 = 1'b0;
  assign po109 = 1'b0;
  assign po110 = 1'b0;
  assign po111 = 1'b0;
  assign po112 = 1'b0;
  assign po113 = 1'b0;
  assign po148 = 1'b0;
  assign po150 = 1'b0;
  assign po012 = po011;
  assign po064 = po051;
  assign po093 = po092;
  assign po121 = po072;
  assign po135 = po134;
  assign po136 = po134;
  assign po137 = po134;
  assign po149 = po002;
endmodule


