// Benchmark "trans_arith" written by ABC on Wed Apr 26 18:25:57 2017

module trans_arith ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119;
  wire n199, n200, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1011, n1012, n1013, n1015, n1016,
    n1017, n1018, n1019, n1021, n1022, n1023, n1024, n1025, n1027, n1028,
    n1029, n1031, n1032, n1033, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1387, n1388, n1390, n1391, n1393,
    n1394, n1396, n1397, n1399, n1400, n1402, n1403, n1405, n1406, n1408,
    n1409, n1411, n1413, n1414, n1416, n1417, n1419, n1420, n1422, n1423,
    n1425, n1426, n1428, n1429, n1431, n1432;
  assign n199 = pi08 & pi24;
  assign n200 = pi73 & n199;
  assign po000 = ~pi75 & n200;
  assign n202 = pi08 & pi25;
  assign n203 = pi09 & pi24;
  assign n204 = ~n202 & ~n203;
  assign n205 = n202 & n203;
  assign n206 = ~n204 & ~n205;
  assign n207 = n200 & n206;
  assign n208 = ~n199 & n204;
  assign n209 = pi73 & ~n208;
  assign n210 = ~pi75 & ~n207;
  assign po001 = n209 & n210;
  assign n212 = pi09 & pi25;
  assign n213 = pi08 & pi26;
  assign n214 = ~n212 & ~n213;
  assign n215 = n212 & n213;
  assign n216 = ~n214 & ~n215;
  assign n217 = pi10 & pi24;
  assign n218 = n216 & n217;
  assign n219 = ~n216 & ~n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = n205 & n220;
  assign n222 = ~n205 & ~n220;
  assign n223 = ~n221 & ~n222;
  assign n224 = pi73 & n223;
  assign n225 = ~n209 & ~n224;
  assign n226 = ~pi75 & ~n225;
  assign n227 = n209 & n223;
  assign po002 = n226 & ~n227;
  assign n229 = ~n218 & ~n221;
  assign n230 = pi09 & pi26;
  assign n231 = pi08 & pi27;
  assign n232 = ~n230 & ~n231;
  assign n233 = n230 & n231;
  assign n234 = ~n232 & ~n233;
  assign n235 = pi10 & pi25;
  assign n236 = n234 & n235;
  assign n237 = ~n234 & ~n235;
  assign n238 = ~n236 & ~n237;
  assign n239 = n215 & n238;
  assign n240 = ~n215 & ~n238;
  assign n241 = ~n239 & ~n240;
  assign n242 = pi11 & pi24;
  assign n243 = n241 & n242;
  assign n244 = ~n241 & ~n242;
  assign n245 = ~n243 & ~n244;
  assign n246 = ~n229 & n245;
  assign n247 = n229 & ~n245;
  assign n248 = ~n246 & ~n247;
  assign n249 = pi73 & n248;
  assign n250 = n225 & ~n249;
  assign n251 = ~pi75 & ~n250;
  assign n252 = n226 & n249;
  assign po003 = n251 & ~n252;
  assign n254 = ~n243 & ~n246;
  assign n255 = ~n236 & ~n239;
  assign n256 = pi09 & pi27;
  assign n257 = pi08 & pi28;
  assign n258 = ~n256 & ~n257;
  assign n259 = n256 & n257;
  assign n260 = ~n258 & ~n259;
  assign n261 = pi10 & pi26;
  assign n262 = n260 & n261;
  assign n263 = ~n260 & ~n261;
  assign n264 = ~n262 & ~n263;
  assign n265 = n233 & n264;
  assign n266 = ~n233 & ~n264;
  assign n267 = ~n265 & ~n266;
  assign n268 = pi11 & pi25;
  assign n269 = n267 & n268;
  assign n270 = ~n267 & ~n268;
  assign n271 = ~n269 & ~n270;
  assign n272 = ~n255 & n271;
  assign n273 = n255 & ~n271;
  assign n274 = ~n272 & ~n273;
  assign n275 = pi12 & pi24;
  assign n276 = n274 & n275;
  assign n277 = ~n274 & ~n275;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~n254 & n278;
  assign n280 = n254 & ~n278;
  assign n281 = ~n279 & ~n280;
  assign n282 = pi73 & n281;
  assign n283 = n250 & ~n282;
  assign n284 = ~pi75 & ~n283;
  assign n285 = n251 & n282;
  assign po004 = n284 & ~n285;
  assign n287 = ~n276 & ~n279;
  assign n288 = ~n269 & ~n272;
  assign n289 = ~n262 & ~n265;
  assign n290 = pi09 & pi28;
  assign n291 = pi08 & pi29;
  assign n292 = ~n290 & ~n291;
  assign n293 = n290 & n291;
  assign n294 = ~n292 & ~n293;
  assign n295 = pi10 & pi27;
  assign n296 = n294 & n295;
  assign n297 = ~n294 & ~n295;
  assign n298 = ~n296 & ~n297;
  assign n299 = n259 & n298;
  assign n300 = ~n259 & ~n298;
  assign n301 = ~n299 & ~n300;
  assign n302 = pi11 & pi26;
  assign n303 = n301 & n302;
  assign n304 = ~n301 & ~n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~n289 & n305;
  assign n307 = n289 & ~n305;
  assign n308 = ~n306 & ~n307;
  assign n309 = pi12 & pi25;
  assign n310 = n308 & n309;
  assign n311 = ~n308 & ~n309;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~n288 & n312;
  assign n314 = n288 & ~n312;
  assign n315 = ~n313 & ~n314;
  assign n316 = pi13 & pi24;
  assign n317 = n315 & n316;
  assign n318 = ~n315 & ~n316;
  assign n319 = ~n317 & ~n318;
  assign n320 = ~n287 & n319;
  assign n321 = n287 & ~n319;
  assign n322 = ~n320 & ~n321;
  assign n323 = pi73 & n322;
  assign n324 = n283 & ~n323;
  assign n325 = n284 & n323;
  assign n326 = ~pi75 & ~n324;
  assign po005 = ~n325 & n326;
  assign n328 = ~n317 & ~n320;
  assign n329 = ~n310 & ~n313;
  assign n330 = ~n303 & ~n306;
  assign n331 = ~n296 & ~n299;
  assign n332 = pi10 & pi28;
  assign n333 = pi09 & pi29;
  assign n334 = pi08 & pi30;
  assign n335 = n333 & ~n334;
  assign n336 = ~n333 & n334;
  assign n337 = ~n335 & ~n336;
  assign n338 = n332 & ~n337;
  assign n339 = ~n332 & n337;
  assign n340 = ~n338 & ~n339;
  assign n341 = n293 & n340;
  assign n342 = ~n293 & ~n340;
  assign n343 = ~n341 & ~n342;
  assign n344 = pi11 & pi27;
  assign n345 = n343 & n344;
  assign n346 = ~n343 & ~n344;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~n331 & n347;
  assign n349 = n331 & ~n347;
  assign n350 = ~n348 & ~n349;
  assign n351 = pi12 & pi26;
  assign n352 = n350 & n351;
  assign n353 = ~n350 & ~n351;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~n330 & n354;
  assign n356 = n330 & ~n354;
  assign n357 = ~n355 & ~n356;
  assign n358 = pi13 & pi25;
  assign n359 = n357 & n358;
  assign n360 = ~n357 & ~n358;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n329 & n361;
  assign n363 = n329 & ~n361;
  assign n364 = ~n362 & ~n363;
  assign n365 = pi14 & pi24;
  assign n366 = n364 & n365;
  assign n367 = ~n364 & ~n365;
  assign n368 = ~n366 & ~n367;
  assign n369 = ~n328 & n368;
  assign n370 = n328 & ~n368;
  assign n371 = ~n369 & ~n370;
  assign n372 = pi73 & n371;
  assign n373 = ~n324 & n372;
  assign n374 = n324 & ~n372;
  assign n375 = ~pi75 & ~n373;
  assign po006 = ~n374 & n375;
  assign n377 = pi11 & pi28;
  assign n378 = ~n366 & ~n369;
  assign n379 = n377 & ~n378;
  assign n380 = ~n377 & n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = pi15 & pi24;
  assign n383 = ~n359 & ~n362;
  assign n384 = n382 & ~n383;
  assign n385 = ~n382 & n383;
  assign n386 = ~n384 & ~n385;
  assign n387 = pi14 & pi25;
  assign n388 = ~n352 & ~n355;
  assign n389 = n387 & ~n388;
  assign n390 = ~n387 & n388;
  assign n391 = ~n389 & ~n390;
  assign n392 = n386 & n391;
  assign n393 = ~n386 & ~n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = pi12 & pi27;
  assign n396 = pi10 & pi29;
  assign n397 = ~n338 & ~n341;
  assign n398 = pi09 & pi30;
  assign n399 = ~n291 & n398;
  assign n400 = n397 & ~n399;
  assign n401 = ~n397 & n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = pi13 & pi26;
  assign n404 = pi08 & pi31;
  assign n405 = ~n345 & ~n348;
  assign n406 = n404 & ~n405;
  assign n407 = ~n404 & n405;
  assign n408 = ~n406 & ~n407;
  assign n409 = n403 & n408;
  assign n410 = ~n403 & ~n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = n402 & ~n411;
  assign n413 = ~n402 & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = n396 & n414;
  assign n416 = ~n396 & ~n414;
  assign n417 = ~n415 & ~n416;
  assign n418 = n395 & ~n417;
  assign n419 = ~n395 & n417;
  assign n420 = ~n418 & ~n419;
  assign n421 = n394 & ~n420;
  assign n422 = ~n394 & n420;
  assign n423 = ~n421 & ~n422;
  assign n424 = n381 & n423;
  assign n425 = ~n381 & ~n423;
  assign n426 = ~n424 & ~n425;
  assign n427 = pi73 & ~n426;
  assign n428 = ~n374 & n427;
  assign n429 = n374 & ~n427;
  assign n430 = ~pi75 & ~n428;
  assign po007 = ~n429 & n430;
  assign n432 = pi72 & pi74;
  assign n433 = ~pi16 & ~pi72;
  assign n434 = pi32 & ~n433;
  assign n435 = ~pi40 & pi72;
  assign n436 = n434 & ~n435;
  assign n437 = ~pi16 & ~pi32;
  assign n438 = ~pi72 & ~n437;
  assign n439 = ~n436 & n438;
  assign n440 = ~n432 & ~n439;
  assign n441 = pi75 & ~n440;
  assign n442 = pi72 & n199;
  assign n443 = ~n200 & ~n442;
  assign n444 = ~pi75 & pi76;
  assign n445 = ~n443 & n444;
  assign po008 = n441 | n445;
  assign n447 = ~pi41 & pi72;
  assign n448 = ~pi17 & ~pi72;
  assign n449 = ~n447 & ~n448;
  assign n450 = pi33 & n449;
  assign n451 = ~pi33 & ~n449;
  assign n452 = ~n450 & ~n451;
  assign n453 = ~n434 & ~n452;
  assign n454 = n436 & n452;
  assign n455 = ~pi72 & ~n453;
  assign n456 = ~n454 & n455;
  assign n457 = ~n432 & ~n456;
  assign n458 = pi75 & ~n457;
  assign n459 = pi73 & n206;
  assign n460 = pi72 & n206;
  assign n461 = ~n459 & ~n460;
  assign n462 = n444 & ~n461;
  assign po009 = n458 | n462;
  assign n464 = ~n450 & ~n454;
  assign n465 = ~pi42 & pi72;
  assign n466 = ~pi18 & ~pi72;
  assign n467 = ~n465 & ~n466;
  assign n468 = pi34 & n467;
  assign n469 = ~pi34 & ~n467;
  assign n470 = ~n468 & ~n469;
  assign n471 = ~n464 & n470;
  assign n472 = n464 & ~n470;
  assign n473 = ~pi72 & ~n471;
  assign n474 = ~n472 & n473;
  assign n475 = ~n432 & ~n474;
  assign n476 = pi75 & ~n475;
  assign n477 = pi72 & n223;
  assign n478 = ~n224 & ~n477;
  assign n479 = n444 & ~n478;
  assign po010 = n476 | n479;
  assign n481 = ~n468 & ~n471;
  assign n482 = ~pi43 & pi72;
  assign n483 = ~pi19 & ~pi72;
  assign n484 = ~n482 & ~n483;
  assign n485 = pi35 & n484;
  assign n486 = ~pi35 & ~n484;
  assign n487 = ~n485 & ~n486;
  assign n488 = ~n481 & n487;
  assign n489 = n481 & ~n487;
  assign n490 = ~pi72 & ~n488;
  assign n491 = ~n489 & n490;
  assign n492 = ~n432 & ~n491;
  assign n493 = pi75 & ~n492;
  assign n494 = pi72 & n248;
  assign n495 = ~n249 & ~n494;
  assign n496 = n444 & ~n495;
  assign po011 = n493 | n496;
  assign n498 = ~n485 & ~n488;
  assign n499 = ~pi44 & pi72;
  assign n500 = ~pi20 & ~pi72;
  assign n501 = ~n499 & ~n500;
  assign n502 = pi36 & n501;
  assign n503 = ~pi36 & ~n501;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~n498 & n504;
  assign n506 = n498 & ~n504;
  assign n507 = ~pi72 & ~n505;
  assign n508 = ~n506 & n507;
  assign n509 = ~n432 & ~n508;
  assign n510 = pi75 & ~n509;
  assign n511 = pi72 & n281;
  assign n512 = ~n282 & ~n511;
  assign n513 = n444 & ~n512;
  assign po012 = n510 | n513;
  assign n515 = ~n502 & ~n505;
  assign n516 = ~pi45 & pi72;
  assign n517 = ~pi21 & ~pi72;
  assign n518 = ~n516 & ~n517;
  assign n519 = pi37 & n518;
  assign n520 = ~pi37 & ~n518;
  assign n521 = ~n519 & ~n520;
  assign n522 = ~n515 & n521;
  assign n523 = n515 & ~n521;
  assign n524 = ~pi72 & ~n522;
  assign n525 = ~n523 & n524;
  assign n526 = ~n432 & ~n525;
  assign n527 = pi75 & ~n526;
  assign n528 = pi72 & n322;
  assign n529 = ~n323 & ~n528;
  assign n530 = n444 & ~n529;
  assign po013 = n527 | n530;
  assign n532 = ~n519 & ~n522;
  assign n533 = ~pi46 & pi72;
  assign n534 = ~pi22 & ~pi72;
  assign n535 = ~n533 & ~n534;
  assign n536 = pi38 & n535;
  assign n537 = ~pi38 & ~n535;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n532 & n538;
  assign n540 = n532 & ~n538;
  assign n541 = ~pi72 & ~n539;
  assign n542 = ~n540 & n541;
  assign n543 = ~n432 & ~n542;
  assign n544 = pi75 & ~n543;
  assign n545 = pi72 & n371;
  assign n546 = ~n372 & ~n545;
  assign n547 = n444 & ~n546;
  assign po014 = n544 | n547;
  assign n549 = ~n536 & ~n539;
  assign n550 = ~pi47 & pi72;
  assign n551 = ~pi23 & ~pi72;
  assign n552 = ~n550 & ~n551;
  assign n553 = pi39 & ~n552;
  assign n554 = ~pi39 & n552;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n549 & ~n555;
  assign n557 = n549 & n555;
  assign n558 = ~pi72 & ~n556;
  assign n559 = ~n557 & n558;
  assign n560 = ~n432 & ~n559;
  assign n561 = pi75 & ~n560;
  assign n562 = pi72 & ~n426;
  assign n563 = ~n427 & ~n562;
  assign n564 = n444 & ~n563;
  assign po015 = n561 | n564;
  assign po048 = pi75 & pi77;
  assign po040 = pi76 & n442;
  assign po016 = po048 | po040;
  assign po041 = pi76 & n460;
  assign po017 = po048 | po041;
  assign po042 = pi76 & n477;
  assign po018 = po048 | po042;
  assign po043 = pi76 & n494;
  assign po019 = po048 | po043;
  assign po044 = pi76 & n511;
  assign po020 = po048 | po044;
  assign po045 = pi76 & n528;
  assign po021 = po048 | po045;
  assign po046 = pi76 & n545;
  assign po022 = po048 | po046;
  assign po047 = pi76 & n562;
  assign po023 = po048 | po047;
  assign n583 = ~pi02 & pi64;
  assign n584 = ~pi04 & pi64;
  assign n585 = pi04 & ~pi64;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~pi66 & ~pi67;
  assign n588 = ~pi68 & ~pi69;
  assign n589 = n587 & n588;
  assign n590 = ~pi70 & ~pi71;
  assign n591 = ~pi65 & n590;
  assign n592 = pi64 & n589;
  assign n593 = n591 & n592;
  assign n594 = pi07 & ~n593;
  assign n595 = ~pi65 & n594;
  assign n596 = ~pi06 & pi64;
  assign n597 = ~n595 & n596;
  assign n598 = pi65 & ~n594;
  assign n599 = ~pi69 & n590;
  assign n600 = ~pi68 & n599;
  assign n601 = ~pi67 & n600;
  assign n602 = ~pi66 & n601;
  assign n603 = ~n598 & n602;
  assign n604 = ~n597 & n603;
  assign n605 = ~pi65 & ~n596;
  assign n606 = n604 & ~n605;
  assign n607 = n594 & ~n606;
  assign n608 = ~pi66 & n607;
  assign n609 = ~pi05 & pi64;
  assign n610 = ~pi65 & ~n609;
  assign n611 = pi65 & n609;
  assign n612 = pi64 & n603;
  assign n613 = pi06 & ~n612;
  assign n614 = n596 & n602;
  assign n615 = n595 & n614;
  assign n616 = ~n613 & ~n615;
  assign n617 = ~n611 & ~n616;
  assign n618 = ~n610 & ~n617;
  assign n619 = ~n608 & n618;
  assign n620 = pi66 & ~n607;
  assign n621 = n601 & ~n620;
  assign n622 = ~n619 & n621;
  assign n623 = n607 & ~n622;
  assign n624 = n608 & ~n618;
  assign n625 = n621 & n624;
  assign n626 = ~n623 & ~n625;
  assign n627 = ~pi67 & ~n626;
  assign n628 = ~n610 & n622;
  assign n629 = ~n611 & n628;
  assign n630 = n616 & ~n629;
  assign n631 = n617 & n628;
  assign n632 = ~n630 & ~n631;
  assign n633 = pi66 & ~n632;
  assign n634 = ~pi66 & n632;
  assign n635 = pi05 & ~pi64;
  assign n636 = ~n609 & ~n635;
  assign n637 = n622 & ~n636;
  assign n638 = pi05 & ~n622;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~pi65 & ~n639;
  assign n641 = pi65 & n639;
  assign n642 = ~n584 & ~n641;
  assign n643 = ~n640 & ~n642;
  assign n644 = ~n634 & n643;
  assign n645 = ~n633 & ~n644;
  assign n646 = ~n627 & ~n645;
  assign n647 = pi67 & n626;
  assign n648 = n600 & ~n647;
  assign n649 = ~n646 & n648;
  assign n650 = ~n640 & n642;
  assign n651 = ~n627 & ~n647;
  assign n652 = ~n633 & ~n634;
  assign n653 = ~n585 & n600;
  assign n654 = n651 & n653;
  assign n655 = n650 & n654;
  assign n656 = n652 & n655;
  assign n657 = ~n649 & ~n656;
  assign n658 = ~n586 & ~n657;
  assign n659 = pi04 & n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n640 & ~n641;
  assign n662 = n584 & ~n661;
  assign n663 = ~n650 & ~n662;
  assign n664 = ~n657 & ~n663;
  assign n665 = n639 & n657;
  assign n666 = ~n664 & ~n665;
  assign n667 = ~pi66 & n666;
  assign n668 = ~pi65 & ~n660;
  assign n669 = pi65 & n660;
  assign n670 = ~pi03 & pi64;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n668 & ~n671;
  assign n673 = ~n667 & n672;
  assign n674 = pi66 & ~n666;
  assign n675 = n632 & n657;
  assign n676 = ~n643 & n652;
  assign n677 = n643 & ~n652;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~n657 & n678;
  assign n680 = ~n675 & ~n679;
  assign n681 = pi67 & n680;
  assign n682 = ~n674 & ~n681;
  assign n683 = ~n673 & n682;
  assign n684 = ~n645 & ~n651;
  assign n685 = n645 & n651;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~n657 & ~n686;
  assign n688 = n626 & n657;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~pi68 & n689;
  assign n691 = ~pi67 & ~n680;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~n683 & n692;
  assign n694 = pi68 & ~n689;
  assign n695 = n599 & ~n694;
  assign n696 = ~n693 & n695;
  assign n697 = ~n660 & ~n696;
  assign n698 = ~n668 & ~n669;
  assign n699 = n670 & ~n698;
  assign n700 = ~n670 & n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = n696 & n701;
  assign n703 = ~n697 & ~n702;
  assign n704 = pi66 & n703;
  assign n705 = ~pi66 & ~n703;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n689 & ~n696;
  assign n708 = ~n690 & ~n694;
  assign n709 = ~n683 & ~n691;
  assign n710 = ~n708 & ~n709;
  assign n711 = n696 & ~n710;
  assign n712 = ~n707 & ~n711;
  assign n713 = pi69 & ~n712;
  assign n714 = ~pi69 & n712;
  assign n715 = ~n713 & ~n714;
  assign n716 = ~n673 & ~n674;
  assign n717 = ~n681 & ~n691;
  assign n718 = ~n716 & ~n717;
  assign n719 = n716 & n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = n696 & ~n720;
  assign n722 = n680 & ~n696;
  assign n723 = ~n721 & ~n722;
  assign n724 = pi68 & ~n723;
  assign n725 = ~pi68 & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = pi03 & ~pi64;
  assign n728 = ~n670 & ~n727;
  assign n729 = n696 & ~n728;
  assign n730 = pi03 & ~n696;
  assign n731 = ~n729 & ~n730;
  assign n732 = pi65 & n731;
  assign n733 = ~pi65 & ~n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n667 & ~n674;
  assign n736 = ~n672 & ~n735;
  assign n737 = n672 & n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = n696 & ~n738;
  assign n740 = n666 & ~n696;
  assign n741 = ~n739 & ~n740;
  assign n742 = pi67 & n741;
  assign n743 = ~pi67 & ~n741;
  assign n744 = ~n742 & ~n743;
  assign n745 = n590 & n706;
  assign n746 = n715 & n726;
  assign n747 = n734 & n744;
  assign n748 = n746 & n747;
  assign n749 = n745 & n748;
  assign n750 = n583 & n749;
  assign n751 = pi02 & ~pi64;
  assign n752 = n749 & ~n751;
  assign n753 = ~n704 & ~n732;
  assign n754 = ~n705 & ~n743;
  assign n755 = ~n753 & n754;
  assign n756 = ~n724 & ~n742;
  assign n757 = ~n755 & n756;
  assign n758 = ~n714 & ~n725;
  assign n759 = ~n757 & n758;
  assign n760 = n590 & ~n713;
  assign n761 = ~n759 & n760;
  assign n762 = ~n752 & ~n761;
  assign n763 = ~n750 & ~n762;
  assign n764 = ~n583 & ~n751;
  assign n765 = n763 & ~n764;
  assign n766 = pi02 & n762;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~pi65 & ~n767;
  assign n769 = ~n583 & ~n734;
  assign n770 = n583 & n734;
  assign n771 = ~n769 & ~n770;
  assign n772 = n763 & ~n771;
  assign n773 = ~n731 & ~n763;
  assign n774 = ~n772 & ~n773;
  assign n775 = pi66 & n774;
  assign n776 = ~pi66 & ~n774;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~n741 & ~n763;
  assign n779 = ~n583 & ~n732;
  assign n780 = ~n733 & ~n779;
  assign n781 = ~n704 & ~n780;
  assign n782 = ~n705 & ~n781;
  assign n783 = n744 & ~n782;
  assign n784 = ~n744 & n782;
  assign n785 = ~n783 & ~n784;
  assign n786 = n763 & n785;
  assign n787 = ~n778 & ~n786;
  assign n788 = pi68 & n787;
  assign n789 = ~pi68 & ~n787;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n706 & ~n780;
  assign n792 = n706 & n780;
  assign n793 = ~n791 & ~n792;
  assign n794 = n763 & ~n793;
  assign n795 = ~n703 & ~n763;
  assign n796 = ~n794 & ~n795;
  assign n797 = pi67 & n796;
  assign n798 = ~pi67 & ~n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n723 & ~n763;
  assign n801 = ~n743 & n782;
  assign n802 = ~n742 & ~n801;
  assign n803 = n726 & ~n802;
  assign n804 = ~n726 & n802;
  assign n805 = n763 & ~n803;
  assign n806 = ~n804 & n805;
  assign n807 = ~n800 & ~n806;
  assign n808 = ~pi69 & n807;
  assign n809 = pi69 & ~n807;
  assign n810 = ~n808 & ~n809;
  assign n811 = n777 & n790;
  assign n812 = n799 & n811;
  assign n813 = n810 & n812;
  assign n814 = ~n768 & n813;
  assign n815 = ~n775 & ~n797;
  assign n816 = ~n789 & ~n798;
  assign n817 = ~n815 & n816;
  assign n818 = ~n788 & ~n809;
  assign n819 = ~n817 & n818;
  assign n820 = ~n808 & ~n819;
  assign n821 = ~n814 & ~n820;
  assign n822 = ~n712 & ~n763;
  assign n823 = ~n724 & n802;
  assign n824 = ~n725 & ~n823;
  assign n825 = ~n715 & ~n824;
  assign n826 = n715 & n824;
  assign n827 = n763 & ~n825;
  assign n828 = ~n826 & n827;
  assign n829 = ~n822 & ~n828;
  assign n830 = ~pi70 & n829;
  assign n831 = ~pi01 & pi64;
  assign n832 = pi65 & n767;
  assign n833 = ~n768 & ~n832;
  assign n834 = ~n831 & n833;
  assign n835 = n813 & n834;
  assign n836 = ~n830 & ~n835;
  assign n837 = ~n821 & n836;
  assign n838 = pi70 & ~n829;
  assign n839 = ~pi71 & ~n838;
  assign n840 = ~n837 & n839;
  assign n841 = pi64 & n840;
  assign n842 = pi01 & ~n841;
  assign n843 = n831 & n840;
  assign n844 = ~n842 & ~n843;
  assign n845 = pi65 & n844;
  assign n846 = ~pi65 & ~n844;
  assign n847 = n767 & ~n840;
  assign n848 = n831 & ~n833;
  assign n849 = ~n834 & ~n848;
  assign n850 = n840 & ~n849;
  assign n851 = ~n847 & ~n850;
  assign n852 = ~pi66 & n851;
  assign n853 = pi66 & ~n851;
  assign n854 = ~pi00 & pi64;
  assign n855 = ~n852 & n854;
  assign n856 = ~n853 & n855;
  assign n857 = ~n845 & ~n846;
  assign n858 = n856 & n857;
  assign n859 = n845 & ~n852;
  assign n860 = ~n853 & ~n859;
  assign n861 = ~n858 & n860;
  assign n862 = ~n831 & ~n832;
  assign n863 = ~n768 & ~n862;
  assign n864 = ~n775 & ~n863;
  assign n865 = ~n776 & ~n864;
  assign n866 = ~n797 & ~n865;
  assign n867 = ~n798 & ~n866;
  assign n868 = ~n790 & ~n867;
  assign n869 = n790 & n867;
  assign n870 = ~n868 & ~n869;
  assign n871 = n840 & ~n870;
  assign n872 = ~n787 & ~n840;
  assign n873 = ~n871 & ~n872;
  assign n874 = pi69 & n873;
  assign n875 = ~n799 & ~n865;
  assign n876 = n799 & n865;
  assign n877 = ~n875 & ~n876;
  assign n878 = n840 & ~n877;
  assign n879 = ~n796 & ~n840;
  assign n880 = ~n878 & ~n879;
  assign n881 = pi68 & n880;
  assign n882 = ~n777 & ~n863;
  assign n883 = n777 & n863;
  assign n884 = ~n882 & ~n883;
  assign n885 = n840 & ~n884;
  assign n886 = ~n774 & ~n840;
  assign n887 = ~n885 & ~n886;
  assign n888 = pi67 & n887;
  assign n889 = ~n881 & ~n888;
  assign n890 = ~pi69 & ~n873;
  assign n891 = ~pi68 & ~n880;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~pi67 & ~n887;
  assign n894 = ~n874 & ~n893;
  assign n895 = n889 & n894;
  assign n896 = n892 & n895;
  assign n897 = ~n861 & n896;
  assign n898 = ~n889 & n892;
  assign n899 = n807 & ~n840;
  assign n900 = ~n789 & n867;
  assign n901 = ~n788 & ~n900;
  assign n902 = ~n810 & ~n901;
  assign n903 = n810 & n901;
  assign n904 = n840 & ~n902;
  assign n905 = ~n903 & n904;
  assign n906 = ~n899 & ~n905;
  assign n907 = pi70 & n906;
  assign n908 = ~n874 & ~n898;
  assign n909 = ~n907 & n908;
  assign n910 = ~n897 & n909;
  assign n911 = ~n829 & ~n840;
  assign n912 = ~n830 & ~n838;
  assign n913 = ~n808 & ~n901;
  assign n914 = ~n809 & ~n913;
  assign n915 = n912 & ~n914;
  assign n916 = ~n912 & n914;
  assign n917 = n840 & ~n915;
  assign n918 = ~n916 & n917;
  assign n919 = ~n911 & ~n918;
  assign n920 = ~pi71 & n919;
  assign n921 = ~pi70 & ~n906;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n910 & n922;
  assign n924 = pi71 & ~n919;
  assign n925 = ~pi64 & n589;
  assign n926 = n591 & n925;
  assign n927 = ~n924 & ~n926;
  assign n928 = ~n923 & n927;
  assign n929 = pi72 & ~n928;
  assign n930 = ~pi72 & n928;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~pi76 & ~n931;
  assign n933 = pi76 & n931;
  assign po064 = n932 | n933;
  assign n935 = n840 & ~n926;
  assign n936 = ~n929 & n935;
  assign n937 = n929 & ~n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~pi76 & ~n938;
  assign n940 = pi76 & n938;
  assign n941 = ~n932 & ~n939;
  assign n942 = ~n940 & n941;
  assign n943 = ~n931 & n939;
  assign po065 = ~n942 & ~n943;
  assign n945 = ~n940 & ~n942;
  assign n946 = n763 & ~n926;
  assign n947 = n937 & ~n946;
  assign n948 = ~n937 & n946;
  assign n949 = ~n947 & ~n948;
  assign n950 = pi76 & n949;
  assign n951 = ~pi76 & ~n949;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n945 & n952;
  assign n954 = n945 & ~n952;
  assign po066 = ~n953 & ~n954;
  assign n956 = ~n950 & ~n953;
  assign n957 = n696 & ~n926;
  assign n958 = ~n947 & n957;
  assign n959 = n947 & ~n957;
  assign n960 = ~n958 & ~n959;
  assign n961 = pi76 & n960;
  assign n962 = ~pi76 & ~n960;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~n956 & n963;
  assign n965 = n956 & ~n963;
  assign po067 = ~n964 & ~n965;
  assign n967 = ~n961 & ~n964;
  assign n968 = ~n657 & ~n926;
  assign n969 = ~n959 & n968;
  assign n970 = n959 & ~n968;
  assign n971 = ~n969 & ~n970;
  assign n972 = pi76 & n971;
  assign n973 = ~pi76 & ~n971;
  assign n974 = ~n972 & ~n973;
  assign n975 = ~n967 & n974;
  assign n976 = n967 & ~n974;
  assign po068 = ~n975 & ~n976;
  assign n978 = ~n972 & ~n975;
  assign n979 = n622 & ~n926;
  assign n980 = ~n970 & n979;
  assign n981 = n970 & ~n979;
  assign n982 = ~n980 & ~n981;
  assign n983 = pi76 & n982;
  assign n984 = ~pi76 & ~n982;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~n978 & n985;
  assign n987 = n978 & ~n985;
  assign po069 = ~n986 & ~n987;
  assign n989 = ~n983 & ~n986;
  assign n990 = n604 & ~n926;
  assign n991 = ~n981 & n990;
  assign n992 = n981 & ~n990;
  assign n993 = ~n991 & ~n992;
  assign n994 = pi76 & n993;
  assign n995 = ~pi76 & ~n993;
  assign n996 = ~n994 & ~n995;
  assign n997 = ~n989 & n996;
  assign n998 = n989 & ~n996;
  assign po070 = ~n997 & ~n998;
  assign n1000 = ~n994 & ~n997;
  assign n1001 = pi07 & n593;
  assign n1002 = pi76 & ~n1001;
  assign n1003 = ~pi76 & n1001;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = n992 & ~n1004;
  assign n1006 = ~n992 & n1004;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = n1000 & n1007;
  assign n1009 = ~n1000 & ~n1007;
  assign po071 = ~n1008 & ~n1009;
  assign n1011 = pi74 & n442;
  assign n1012 = pi73 & ~n1011;
  assign n1013 = ~pi73 & n1011;
  assign po080 = n1012 | n1013;
  assign n1015 = ~n208 & n432;
  assign n1016 = pi73 & ~n1015;
  assign n1017 = n206 & n1011;
  assign n1018 = ~n1012 & n1015;
  assign n1019 = ~n1017 & n1018;
  assign po081 = n1016 | n1019;
  assign n1021 = ~pi73 & n208;
  assign n1022 = pi74 & n477;
  assign n1023 = ~n1021 & n1022;
  assign n1024 = ~n1015 & ~n1022;
  assign n1025 = ~pi73 & n1024;
  assign po082 = ~n1023 & ~n1025;
  assign n1027 = pi74 & n494;
  assign n1028 = ~n1025 & n1027;
  assign n1029 = n1025 & ~n1027;
  assign po083 = ~n1028 & ~n1029;
  assign n1031 = pi74 & n511;
  assign n1032 = ~n1029 & n1031;
  assign n1033 = n1029 & ~n1031;
  assign po084 = ~n1032 & ~n1033;
  assign n1035 = n1024 & ~n1027;
  assign n1036 = ~n1031 & n1035;
  assign n1037 = pi74 & n528;
  assign n1038 = n1036 & ~n1037;
  assign n1039 = n1016 & n1038;
  assign n1040 = ~n1036 & n1037;
  assign n1041 = ~n1038 & ~n1040;
  assign n1042 = n1016 & n1037;
  assign n1043 = n1041 & ~n1042;
  assign po085 = n1039 | n1043;
  assign n1045 = pi74 & n545;
  assign n1046 = n1041 & n1045;
  assign n1047 = ~n1041 & ~n1045;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1040 & ~n1048;
  assign n1050 = n545 & n1040;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = n1039 & ~n1051;
  assign n1053 = ~n1039 & n1051;
  assign po086 = n1052 | n1053;
  assign n1055 = ~n1039 & n1049;
  assign n1056 = n432 & ~n1046;
  assign n1057 = ~n426 & n1056;
  assign n1058 = n426 & n1046;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = n1055 & ~n1059;
  assign n1061 = ~n1055 & n1059;
  assign po087 = n1060 | n1061;
  assign n1063 = pi75 & n442;
  assign n1064 = ~pi48 & pi56;
  assign n1065 = pi48 & ~pi56;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = pi72 & ~n1066;
  assign n1068 = ~n1063 & n1067;
  assign n1069 = n1063 & n1066;
  assign po088 = n1068 | n1069;
  assign n1071 = pi75 & n460;
  assign n1072 = pi74 & n206;
  assign n1073 = n1067 & n1072;
  assign n1074 = pi74 & n199;
  assign n1075 = ~n1067 & ~n1074;
  assign n1076 = pi49 & ~pi57;
  assign n1077 = ~pi49 & pi57;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n1064 & ~n1078;
  assign n1080 = ~n1064 & n1078;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = pi72 & n1081;
  assign n1083 = ~n1075 & n1082;
  assign n1084 = ~n1073 & ~n1083;
  assign n1085 = n1067 & n1081;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = n1071 & ~n1086;
  assign n1088 = ~n1071 & n1086;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n1068 & n1089;
  assign n1091 = n1068 & ~n1089;
  assign po089 = ~n1090 & ~n1091;
  assign n1093 = ~n1087 & ~n1090;
  assign n1094 = pi75 & n477;
  assign n1095 = pi72 & ~n1075;
  assign n1096 = ~n1076 & ~n1080;
  assign n1097 = pi50 & ~pi58;
  assign n1098 = ~pi50 & pi58;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = ~n1096 & n1099;
  assign n1101 = n1096 & ~n1099;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = n1095 & n1102;
  assign n1104 = ~n1082 & ~n1103;
  assign n1105 = n1082 & n1103;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = pi74 & n223;
  assign n1108 = pi72 & n1102;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = n1067 & ~n1109;
  assign n1111 = n1106 & n1110;
  assign n1112 = ~n1106 & ~n1110;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = n1085 & n1113;
  assign n1115 = ~n1085 & ~n1113;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = n1094 & ~n1116;
  assign n1118 = ~n1094 & n1116;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1093 & n1119;
  assign n1121 = n1093 & ~n1119;
  assign po090 = ~n1120 & ~n1121;
  assign n1123 = ~n1117 & ~n1120;
  assign n1124 = pi75 & n494;
  assign n1125 = ~n1111 & ~n1114;
  assign n1126 = ~n1072 & ~n1082;
  assign n1127 = n1108 & ~n1126;
  assign n1128 = ~n1097 & ~n1100;
  assign n1129 = pi51 & ~pi59;
  assign n1130 = ~pi51 & pi59;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = n1128 & ~n1131;
  assign n1133 = ~n1128 & n1131;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = n1095 & n1134;
  assign n1136 = ~n1127 & ~n1135;
  assign n1137 = pi72 & n1134;
  assign n1138 = ~n1126 & n1137;
  assign n1139 = n1103 & n1138;
  assign n1140 = ~n1136 & ~n1139;
  assign n1141 = n1082 & ~n1109;
  assign n1142 = n1140 & n1141;
  assign n1143 = ~n1140 & ~n1141;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = n1105 & n1144;
  assign n1146 = ~n1105 & ~n1144;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = pi74 & n248;
  assign n1149 = ~n1137 & ~n1148;
  assign n1150 = n1067 & ~n1149;
  assign n1151 = n1147 & n1150;
  assign n1152 = ~n1147 & ~n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1125 & n1153;
  assign n1155 = n1125 & ~n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = n1124 & ~n1156;
  assign n1158 = ~n1124 & n1156;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = ~n1123 & n1159;
  assign n1161 = n1123 & ~n1159;
  assign po091 = ~n1160 & ~n1161;
  assign n1163 = ~n1157 & ~n1160;
  assign n1164 = pi75 & n511;
  assign n1165 = ~n1151 & ~n1154;
  assign n1166 = ~n1142 & ~n1145;
  assign n1167 = n1082 & ~n1149;
  assign n1168 = ~n1129 & ~n1133;
  assign n1169 = pi52 & ~pi60;
  assign n1170 = ~pi52 & pi60;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = n1168 & ~n1171;
  assign n1173 = ~n1168 & n1171;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = n1095 & n1174;
  assign n1176 = ~n1138 & ~n1175;
  assign n1177 = n1108 & n1176;
  assign n1178 = ~n1108 & ~n1176;
  assign n1179 = ~n1139 & ~n1178;
  assign n1180 = pi72 & n1174;
  assign n1181 = ~n1126 & n1180;
  assign n1182 = n1135 & n1181;
  assign n1183 = ~n1179 & ~n1182;
  assign n1184 = ~n1177 & ~n1183;
  assign n1185 = n1167 & ~n1184;
  assign n1186 = ~n1167 & n1184;
  assign n1187 = ~n1185 & ~n1186;
  assign n1188 = ~n1166 & n1187;
  assign n1189 = n1166 & ~n1187;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = pi74 & n281;
  assign n1192 = ~n1180 & ~n1191;
  assign n1193 = n1067 & ~n1192;
  assign n1194 = n1190 & n1193;
  assign n1195 = ~n1190 & ~n1193;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1165 & n1196;
  assign n1198 = n1165 & ~n1196;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = n1164 & ~n1199;
  assign n1201 = ~n1164 & n1199;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1163 & n1202;
  assign n1204 = n1163 & ~n1202;
  assign po092 = ~n1203 & ~n1204;
  assign n1206 = ~n1200 & ~n1203;
  assign n1207 = pi75 & n528;
  assign n1208 = ~n1194 & ~n1197;
  assign n1209 = ~n1185 & ~n1188;
  assign n1210 = ~n1169 & ~n1173;
  assign n1211 = pi53 & ~pi61;
  assign n1212 = ~pi53 & pi61;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = n1210 & ~n1213;
  assign n1215 = ~n1210 & n1213;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = n1095 & n1216;
  assign n1218 = ~n1181 & ~n1217;
  assign n1219 = pi72 & n1216;
  assign n1220 = ~n1126 & n1219;
  assign n1221 = n1175 & n1220;
  assign n1222 = ~n1218 & ~n1221;
  assign n1223 = ~n1109 & n1137;
  assign n1224 = n1222 & n1223;
  assign n1225 = ~n1222 & ~n1223;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = n1182 & n1226;
  assign n1228 = ~n1182 & ~n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = n1108 & ~n1149;
  assign n1231 = n1229 & n1230;
  assign n1232 = ~n1229 & ~n1230;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = n1108 & ~n1176;
  assign n1235 = n1233 & n1234;
  assign n1236 = ~n1233 & ~n1234;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = n1082 & ~n1192;
  assign n1239 = n1237 & n1238;
  assign n1240 = ~n1237 & ~n1238;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = ~n1209 & n1241;
  assign n1243 = n1209 & ~n1241;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = pi74 & n322;
  assign n1246 = ~n1219 & ~n1245;
  assign n1247 = n1067 & ~n1246;
  assign n1248 = n1244 & n1247;
  assign n1249 = ~n1244 & ~n1247;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~n1208 & n1250;
  assign n1252 = n1208 & ~n1250;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = n1207 & ~n1253;
  assign n1255 = ~n1207 & n1253;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n1206 & n1256;
  assign n1258 = n1206 & ~n1256;
  assign po093 = ~n1257 & ~n1258;
  assign n1260 = ~n1254 & ~n1257;
  assign n1261 = pi75 & n545;
  assign n1262 = ~n1248 & ~n1251;
  assign n1263 = ~n1239 & ~n1242;
  assign n1264 = ~n1231 & ~n1235;
  assign n1265 = ~n1224 & ~n1227;
  assign n1266 = ~n1109 & n1180;
  assign n1267 = ~n1211 & ~n1215;
  assign n1268 = pi54 & ~pi62;
  assign n1269 = ~pi54 & pi62;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1267 & n1270;
  assign n1272 = n1267 & ~n1270;
  assign n1273 = pi72 & ~n1271;
  assign n1274 = ~n1272 & n1273;
  assign n1275 = ~n1075 & n1274;
  assign n1276 = ~n1220 & n1275;
  assign n1277 = n1220 & ~n1275;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = n1266 & ~n1278;
  assign n1280 = ~n1266 & n1278;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = n1221 & n1281;
  assign n1283 = ~n1221 & ~n1281;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = n1137 & n1284;
  assign n1286 = ~n1137 & ~n1284;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = ~n1265 & n1287;
  assign n1289 = n1265 & ~n1287;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = n1108 & ~n1192;
  assign n1292 = n1290 & n1291;
  assign n1293 = ~n1290 & ~n1291;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n1264 & n1294;
  assign n1296 = n1264 & ~n1294;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = n1082 & ~n1246;
  assign n1299 = n1297 & n1298;
  assign n1300 = ~n1297 & ~n1298;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = ~n1263 & n1301;
  assign n1303 = n1263 & ~n1301;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = pi74 & n371;
  assign n1306 = ~n1274 & ~n1305;
  assign n1307 = n1067 & ~n1306;
  assign n1308 = n1304 & n1307;
  assign n1309 = ~n1304 & ~n1307;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1262 & n1310;
  assign n1312 = n1262 & ~n1310;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = n1261 & ~n1313;
  assign n1315 = ~n1261 & n1313;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = ~n1260 & n1316;
  assign n1318 = n1260 & ~n1316;
  assign po094 = ~n1317 & ~n1318;
  assign n1320 = ~n1285 & ~n1288;
  assign n1321 = n1108 & n1216;
  assign n1322 = ~n1108 & ~n1219;
  assign n1323 = ~n1109 & ~n1321;
  assign n1324 = ~n1322 & n1323;
  assign n1325 = ~n1246 & n1324;
  assign n1326 = n1320 & ~n1325;
  assign n1327 = ~n1320 & n1325;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1126 & ~n1217;
  assign n1330 = n1274 & n1329;
  assign n1331 = ~n1134 & n1174;
  assign n1332 = n1027 & n1331;
  assign n1333 = n1134 & ~n1174;
  assign n1334 = n1031 & n1333;
  assign n1335 = ~n1332 & ~n1334;
  assign n1336 = n1330 & ~n1335;
  assign n1337 = ~n1330 & n1335;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~n1292 & ~n1295;
  assign n1340 = n1082 & ~n1306;
  assign n1341 = ~n1268 & ~n1271;
  assign n1342 = ~pi55 & ~pi63;
  assign n1343 = pi55 & pi63;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = n1341 & ~n1344;
  assign n1346 = ~n1341 & n1344;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = n1095 & ~n1347;
  assign n1349 = n1340 & ~n1348;
  assign n1350 = ~n1340 & n1348;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = n1339 & n1351;
  assign n1353 = ~n1339 & ~n1351;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = n1338 & ~n1354;
  assign n1356 = ~n1338 & n1354;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = pi75 & n562;
  assign n1359 = ~n1314 & ~n1317;
  assign n1360 = n1358 & ~n1359;
  assign n1361 = ~n1358 & n1359;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1299 & ~n1302;
  assign n1364 = n1362 & ~n1363;
  assign n1365 = ~n1362 & n1363;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = n1357 & n1366;
  assign n1368 = ~n1357 & ~n1366;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = ~n1308 & ~n1311;
  assign n1371 = ~n1279 & ~n1282;
  assign n1372 = n1370 & ~n1371;
  assign n1373 = ~n1370 & n1371;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = pi74 & ~n426;
  assign n1376 = n1347 & ~n1375;
  assign n1377 = n1067 & ~n1376;
  assign n1378 = n1374 & ~n1377;
  assign n1379 = ~n1374 & n1377;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = n1369 & ~n1380;
  assign n1382 = ~n1369 & n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = n1328 & n1383;
  assign n1385 = ~n1328 & ~n1383;
  assign po095 = n1384 | n1385;
  assign n1387 = pi73 & n440;
  assign n1388 = ~pi73 & ~n440;
  assign po104 = n1387 | n1388;
  assign n1390 = ~n456 & n1387;
  assign n1391 = ~n457 & ~n1387;
  assign po105 = n1390 | n1391;
  assign n1393 = n475 & n1390;
  assign n1394 = ~n475 & ~n1390;
  assign po106 = n1393 | n1394;
  assign n1396 = ~n491 & n1393;
  assign n1397 = ~n492 & ~n1393;
  assign po107 = n1396 | n1397;
  assign n1399 = n509 & n1396;
  assign n1400 = ~n509 & ~n1396;
  assign po108 = n1399 | n1400;
  assign n1402 = ~n526 & ~n1399;
  assign n1403 = ~n525 & n1399;
  assign po109 = n1402 | n1403;
  assign n1405 = n543 & n1403;
  assign n1406 = ~n543 & ~n1403;
  assign po110 = n1405 | n1406;
  assign n1408 = ~n559 & n1405;
  assign n1409 = ~n560 & ~n1405;
  assign po111 = n1408 | n1409;
  assign n1411 = pi75 & ~n200;
  assign po112 = po000 | n1411;
  assign n1413 = n459 & ~n1411;
  assign n1414 = pi75 & ~n209;
  assign po113 = n1413 | n1414;
  assign n1416 = n224 & ~n1414;
  assign n1417 = pi75 & n225;
  assign po114 = n1416 | n1417;
  assign n1419 = n249 & ~n1417;
  assign n1420 = ~n249 & n1417;
  assign po115 = n1419 | n1420;
  assign n1422 = n282 & ~n1420;
  assign n1423 = pi75 & n283;
  assign po116 = n1422 | n1423;
  assign n1425 = n323 & ~n1423;
  assign n1426 = ~n323 & n1423;
  assign po117 = n1425 | n1426;
  assign n1428 = n372 & ~n1426;
  assign n1429 = pi75 & n374;
  assign po118 = n1428 | n1429;
  assign n1431 = n427 & ~n1429;
  assign n1432 = ~n427 & n1429;
  assign po119 = n1431 | n1432;
  assign po024 = pi72;
  assign po025 = pi72;
  assign po026 = pi72;
  assign po027 = pi72;
  assign po028 = pi72;
  assign po029 = pi72;
  assign po030 = pi72;
  assign po031 = pi72;
  assign po032 = pi77;
  assign po033 = pi77;
  assign po034 = pi77;
  assign po035 = pi77;
  assign po036 = pi77;
  assign po037 = pi77;
  assign po038 = pi77;
  assign po039 = pi77;
  assign po049 = po048;
  assign po050 = po048;
  assign po051 = po048;
  assign po052 = po048;
  assign po053 = po048;
  assign po054 = po048;
  assign po055 = po048;
  assign po056 = po016;
  assign po057 = po017;
  assign po058 = po018;
  assign po059 = po019;
  assign po060 = po020;
  assign po061 = po021;
  assign po062 = po022;
  assign po063 = po023;
  assign po072 = po064;
  assign po073 = po065;
  assign po074 = po066;
  assign po075 = po067;
  assign po076 = po068;
  assign po077 = po069;
  assign po078 = po070;
  assign po079 = po071;
  assign po096 = po088;
  assign po097 = po089;
  assign po098 = po090;
  assign po099 = po091;
  assign po100 = po092;
  assign po101 = po093;
  assign po102 = po094;
  assign po103 = po095;
endmodule


