// Benchmark "top" written by ABC on Wed Apr 26 18:13:28 2017

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
    n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
    n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
    n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
    n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
    n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
    n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
    n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
    n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
    n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
    n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
    n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
    n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
    n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
    n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
    n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
    n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
    n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
    n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
    n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
    n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
    n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
    n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
    n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
    n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
    n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
    n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
    n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
    n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
    n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
    n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
    n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
    n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
    n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
    n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
    n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
    n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
    n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
    n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
    n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
    n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
    n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
    n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
    n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
    n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
    n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
    n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
    n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
    n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
    n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
    n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
    n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
    n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
    n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
    n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
    n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
    n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
    n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
    n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
    n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
    n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
    n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
    n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
    n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
    n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
    n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
    n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
    n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
    n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
    n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
    n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
    n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
    n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7062, n7063, n7065;
  assign n65 = ~pi19 & ~pi20;
  assign n66 = ~pi30 & ~pi31;
  assign n67 = ~pi29 & n66;
  assign n68 = ~pi25 & ~pi26;
  assign n69 = ~pi27 & ~pi28;
  assign n70 = n68 & n69;
  assign n71 = n67 & n70;
  assign n72 = ~pi23 & ~pi24;
  assign n73 = n71 & n72;
  assign n74 = ~pi22 & n73;
  assign n75 = ~pi21 & n74;
  assign n76 = n65 & n75;
  assign n77 = ~pi15 & ~pi16;
  assign n78 = ~pi17 & ~pi18;
  assign n79 = n77 & n78;
  assign n80 = n76 & n79;
  assign n81 = ~pi14 & n80;
  assign n82 = ~pi13 & n81;
  assign n83 = ~pi12 & n82;
  assign n84 = ~pi00 & ~pi01;
  assign n85 = ~pi02 & n84;
  assign n86 = ~pi03 & n85;
  assign n87 = ~pi10 & ~pi11;
  assign n88 = ~pi09 & ~pi12;
  assign n89 = n87 & n88;
  assign n90 = n82 & n89;
  assign n91 = ~pi07 & ~pi08;
  assign n92 = n90 & n91;
  assign n93 = ~pi06 & n92;
  assign n94 = ~pi04 & ~pi05;
  assign n95 = n93 & n94;
  assign n96 = pi03 & ~n85;
  assign n97 = ~n86 & ~n96;
  assign n98 = n95 & n97;
  assign n99 = ~pi05 & n93;
  assign n100 = ~pi04 & ~n98;
  assign n101 = ~pi03 & n95;
  assign n102 = pi00 & pi01;
  assign n103 = pi02 & ~n84;
  assign n104 = ~n102 & n103;
  assign n105 = n101 & n104;
  assign n106 = pi02 & ~n105;
  assign n107 = ~pi03 & ~n106;
  assign n108 = ~n100 & ~n107;
  assign n109 = ~pi02 & n102;
  assign n110 = n101 & n109;
  assign n111 = ~n106 & ~n110;
  assign n112 = pi02 & pi03;
  assign n113 = ~n85 & ~n103;
  assign n114 = ~n112 & ~n113;
  assign n115 = n95 & n114;
  assign n116 = pi00 & n115;
  assign n117 = ~pi01 & n116;
  assign n118 = ~pi03 & n99;
  assign n119 = ~n100 & n118;
  assign n120 = ~n117 & n119;
  assign n121 = n111 & n120;
  assign n122 = n99 & ~n108;
  assign n123 = ~n121 & n122;
  assign n124 = n84 & n119;
  assign n125 = n111 & n124;
  assign n126 = ~n123 & ~n125;
  assign n127 = ~n84 & ~n117;
  assign n128 = ~n110 & n127;
  assign n129 = n107 & ~n128;
  assign n130 = pi04 & ~n129;
  assign n131 = ~pi04 & n129;
  assign n132 = ~n130 & ~n131;
  assign n133 = ~n126 & n132;
  assign n134 = ~n98 & n133;
  assign n135 = n98 & ~n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = ~pi05 & n136;
  assign n138 = pi05 & ~n136;
  assign n139 = ~n137 & ~n138;
  assign n140 = ~pi00 & ~n126;
  assign n141 = ~n116 & ~n140;
  assign n142 = ~pi01 & ~n126;
  assign n143 = ~n141 & ~n142;
  assign n144 = pi00 & ~n126;
  assign n145 = ~pi01 & n144;
  assign n146 = ~n115 & n145;
  assign n147 = ~n143 & ~n146;
  assign n148 = ~pi02 & ~n147;
  assign n149 = ~n105 & ~n110;
  assign n150 = n126 & ~n149;
  assign n151 = n111 & ~n127;
  assign n152 = ~n111 & n127;
  assign n153 = ~n151 & ~n152;
  assign n154 = ~n126 & n153;
  assign n155 = ~n150 & ~n154;
  assign n156 = ~pi03 & ~n155;
  assign n157 = pi02 & ~n141;
  assign n158 = n145 & ~n157;
  assign n159 = ~n156 & ~n158;
  assign n160 = ~n148 & n159;
  assign n161 = ~n96 & ~n129;
  assign n162 = ~n126 & n161;
  assign n163 = pi04 & ~n162;
  assign n164 = pi03 & n155;
  assign n165 = ~n163 & ~n164;
  assign n166 = ~n160 & n165;
  assign n167 = ~pi04 & n162;
  assign n168 = ~n137 & ~n167;
  assign n169 = ~n166 & n168;
  assign n170 = n93 & ~n138;
  assign n171 = ~n169 & n170;
  assign n172 = ~n156 & ~n164;
  assign n173 = pi02 & n147;
  assign n174 = ~n163 & ~n167;
  assign n175 = n84 & n92;
  assign n176 = ~pi06 & n175;
  assign n177 = n174 & n176;
  assign n178 = n172 & n177;
  assign n179 = n139 & n178;
  assign n180 = ~n148 & ~n173;
  assign n181 = n179 & n180;
  assign n182 = ~n171 & ~n181;
  assign n183 = ~pi05 & n182;
  assign n184 = ~n84 & ~n145;
  assign n185 = ~n173 & ~n184;
  assign n186 = ~n148 & ~n185;
  assign n187 = ~n164 & ~n186;
  assign n188 = ~n156 & ~n187;
  assign n189 = ~n163 & ~n188;
  assign n190 = ~n167 & ~n189;
  assign n191 = ~n182 & ~n190;
  assign n192 = ~n183 & ~n191;
  assign n193 = n139 & ~n192;
  assign n194 = ~n139 & n192;
  assign n195 = ~n193 & ~n194;
  assign n196 = ~n162 & n182;
  assign n197 = ~n174 & ~n188;
  assign n198 = n174 & n188;
  assign n199 = ~n182 & ~n197;
  assign n200 = ~n198 & n199;
  assign n201 = ~n196 & ~n200;
  assign n202 = ~pi05 & n201;
  assign n203 = ~pi06 & n195;
  assign n204 = ~n172 & ~n186;
  assign n205 = n172 & n186;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n182 & ~n206;
  assign n208 = ~n155 & n182;
  assign n209 = ~n207 & ~n208;
  assign n210 = ~pi04 & ~n209;
  assign n211 = n113 & n141;
  assign n212 = ~n157 & ~n211;
  assign n213 = ~n182 & n212;
  assign n214 = n147 & n182;
  assign n215 = ~n213 & ~n214;
  assign n216 = ~pi03 & n215;
  assign n217 = pi00 & ~n123;
  assign n218 = ~pi01 & ~n217;
  assign n219 = pi01 & n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = ~n182 & ~n220;
  assign n222 = ~n144 & n182;
  assign n223 = ~n221 & ~n222;
  assign n224 = pi02 & ~n223;
  assign n225 = ~n216 & n224;
  assign n226 = pi04 & n209;
  assign n227 = pi03 & ~n215;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n225 & n228;
  assign n230 = ~n210 & ~n229;
  assign n231 = pi05 & ~n201;
  assign n232 = ~pi02 & n223;
  assign n233 = ~n224 & ~n232;
  assign n234 = ~n210 & ~n226;
  assign n235 = ~n216 & ~n227;
  assign n236 = n234 & n235;
  assign n237 = pi00 & ~n182;
  assign n238 = ~pi01 & n237;
  assign n239 = n233 & ~n238;
  assign n240 = n236 & n239;
  assign n241 = ~n230 & ~n231;
  assign n242 = ~n240 & n241;
  assign n243 = ~n202 & ~n203;
  assign n244 = ~n242 & n243;
  assign n245 = pi06 & ~n195;
  assign n246 = n92 & ~n245;
  assign n247 = ~n244 & n246;
  assign n248 = ~n202 & ~n231;
  assign n249 = ~n203 & ~n245;
  assign n250 = n175 & n233;
  assign n251 = n236 & n250;
  assign n252 = n248 & n251;
  assign n253 = n249 & n252;
  assign n254 = ~n247 & ~n253;
  assign n255 = ~n195 & n254;
  assign n256 = ~n84 & ~n238;
  assign n257 = ~n224 & ~n256;
  assign n258 = ~n232 & ~n257;
  assign n259 = ~n216 & n258;
  assign n260 = n228 & ~n259;
  assign n261 = ~n210 & ~n260;
  assign n262 = ~n202 & n261;
  assign n263 = ~n231 & ~n262;
  assign n264 = n249 & ~n263;
  assign n265 = ~n249 & n263;
  assign n266 = ~n254 & ~n264;
  assign n267 = ~n265 & n266;
  assign n268 = ~n255 & ~n267;
  assign n269 = ~pi07 & n268;
  assign n270 = ~n215 & n254;
  assign n271 = ~n235 & ~n258;
  assign n272 = n235 & n258;
  assign n273 = ~n271 & ~n272;
  assign n274 = ~n254 & n273;
  assign n275 = ~n270 & ~n274;
  assign n276 = ~pi04 & n275;
  assign n277 = ~n223 & n254;
  assign n278 = ~n233 & ~n256;
  assign n279 = n233 & n256;
  assign n280 = ~n278 & ~n279;
  assign n281 = ~n254 & n280;
  assign n282 = ~n277 & ~n281;
  assign n283 = pi03 & ~n282;
  assign n284 = ~n276 & n283;
  assign n285 = pi04 & ~n275;
  assign n286 = n209 & n254;
  assign n287 = ~n227 & ~n259;
  assign n288 = n234 & ~n287;
  assign n289 = ~n234 & n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n254 & n290;
  assign n292 = ~n286 & ~n291;
  assign n293 = pi05 & ~n292;
  assign n294 = ~n285 & ~n293;
  assign n295 = ~n284 & n294;
  assign n296 = ~n201 & n254;
  assign n297 = ~n248 & ~n261;
  assign n298 = n248 & n261;
  assign n299 = ~n297 & ~n298;
  assign n300 = ~n254 & n299;
  assign n301 = ~n296 & ~n300;
  assign n302 = ~pi06 & n301;
  assign n303 = ~pi05 & n292;
  assign n304 = ~n302 & ~n303;
  assign n305 = ~n295 & n304;
  assign n306 = pi07 & ~n268;
  assign n307 = pi06 & ~n301;
  assign n308 = ~n306 & ~n307;
  assign n309 = ~n305 & n308;
  assign n310 = ~n269 & ~n309;
  assign n311 = ~pi08 & n90;
  assign n312 = ~n269 & ~n306;
  assign n313 = ~n293 & ~n303;
  assign n314 = ~n84 & ~n102;
  assign n315 = pi00 & n171;
  assign n316 = n314 & ~n315;
  assign n317 = ~n314 & n315;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~n254 & ~n318;
  assign n320 = n237 & n254;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~pi02 & ~n321;
  assign n323 = ~n302 & ~n307;
  assign n324 = ~pi03 & n282;
  assign n325 = ~n283 & ~n324;
  assign n326 = ~n276 & ~n285;
  assign n327 = n311 & ~n322;
  assign n328 = n313 & n327;
  assign n329 = n323 & n325;
  assign n330 = n326 & n329;
  assign n331 = n312 & n328;
  assign n332 = n330 & n331;
  assign n333 = n311 & ~n332;
  assign n334 = ~n310 & n333;
  assign n335 = pi02 & n321;
  assign n336 = n332 & ~n335;
  assign n337 = pi00 & n254;
  assign n338 = ~pi01 & ~n337;
  assign n339 = n336 & n338;
  assign n340 = ~n334 & ~n339;
  assign n341 = ~n268 & n340;
  assign n342 = ~n335 & n338;
  assign n343 = ~n322 & ~n342;
  assign n344 = ~n324 & n343;
  assign n345 = ~n283 & ~n344;
  assign n346 = ~n276 & ~n345;
  assign n347 = ~n285 & ~n346;
  assign n348 = ~n303 & ~n347;
  assign n349 = ~n293 & ~n348;
  assign n350 = ~n302 & ~n349;
  assign n351 = ~n307 & ~n350;
  assign n352 = n312 & ~n351;
  assign n353 = ~n312 & n351;
  assign n354 = ~n340 & ~n352;
  assign n355 = ~n353 & n354;
  assign n356 = ~n341 & ~n355;
  assign n357 = pi08 & ~n356;
  assign n358 = ~pi08 & n356;
  assign n359 = n301 & n340;
  assign n360 = ~n323 & ~n349;
  assign n361 = n323 & n349;
  assign n362 = ~n340 & ~n360;
  assign n363 = ~n361 & n362;
  assign n364 = ~n359 & ~n363;
  assign n365 = pi07 & n364;
  assign n366 = ~n292 & n340;
  assign n367 = n313 & ~n347;
  assign n368 = ~n313 & n347;
  assign n369 = ~n340 & ~n367;
  assign n370 = ~n368 & n369;
  assign n371 = ~n366 & ~n370;
  assign n372 = ~pi06 & n371;
  assign n373 = n282 & n340;
  assign n374 = n325 & ~n343;
  assign n375 = ~n325 & n343;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n340 & n376;
  assign n378 = ~n373 & ~n377;
  assign n379 = pi04 & n378;
  assign n380 = ~n322 & ~n335;
  assign n381 = ~n338 & ~n380;
  assign n382 = n338 & n380;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n340 & ~n383;
  assign n385 = n321 & n340;
  assign n386 = ~n384 & ~n385;
  assign n387 = pi03 & ~n386;
  assign n388 = ~n379 & ~n387;
  assign n389 = ~n326 & ~n345;
  assign n390 = n326 & n345;
  assign n391 = ~n389 & ~n390;
  assign n392 = ~n340 & ~n391;
  assign n393 = ~n275 & n340;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~pi05 & n394;
  assign n396 = ~pi04 & ~n378;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n388 & n397;
  assign n399 = pi05 & ~n394;
  assign n400 = pi06 & ~n371;
  assign n401 = ~n399 & ~n400;
  assign n402 = ~n398 & n401;
  assign n403 = ~n372 & ~n402;
  assign n404 = ~n365 & ~n403;
  assign n405 = ~pi07 & ~n364;
  assign n406 = ~n358 & ~n405;
  assign n407 = ~n404 & n406;
  assign n408 = n90 & ~n357;
  assign n409 = ~n407 & n408;
  assign n410 = ~n357 & ~n358;
  assign n411 = ~n365 & ~n405;
  assign n412 = ~pi03 & n386;
  assign n413 = ~n387 & ~n412;
  assign n414 = ~n395 & ~n399;
  assign n415 = ~n379 & ~n396;
  assign n416 = ~n372 & ~n400;
  assign n417 = n90 & n413;
  assign n418 = n414 & n415;
  assign n419 = n417 & n418;
  assign n420 = n416 & n419;
  assign n421 = n411 & n420;
  assign n422 = n410 & n421;
  assign n423 = ~n409 & ~n422;
  assign n424 = pi00 & n247;
  assign n425 = n314 & ~n424;
  assign n426 = ~n314 & n424;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~n340 & ~n427;
  assign n429 = pi00 & ~n254;
  assign n430 = n340 & n429;
  assign n431 = ~n428 & ~n430;
  assign n432 = pi02 & n431;
  assign n433 = ~pi02 & ~n431;
  assign n434 = pi00 & ~n340;
  assign n435 = ~pi01 & n434;
  assign n436 = ~n433 & ~n435;
  assign n437 = ~n432 & ~n436;
  assign n438 = n422 & ~n437;
  assign n439 = ~n423 & ~n438;
  assign n440 = ~n432 & ~n433;
  assign n441 = n84 & n440;
  assign n442 = n422 & n441;
  assign n443 = ~n439 & ~n442;
  assign n444 = ~n356 & n443;
  assign n445 = ~n84 & ~n435;
  assign n446 = ~n432 & ~n445;
  assign n447 = ~n433 & ~n446;
  assign n448 = ~n387 & ~n447;
  assign n449 = ~n412 & ~n448;
  assign n450 = ~n379 & ~n449;
  assign n451 = ~n396 & ~n450;
  assign n452 = ~n395 & n451;
  assign n453 = ~n399 & ~n452;
  assign n454 = ~n400 & n453;
  assign n455 = ~n372 & ~n454;
  assign n456 = ~n365 & ~n455;
  assign n457 = ~n405 & ~n456;
  assign n458 = ~n410 & ~n457;
  assign n459 = n410 & n457;
  assign n460 = ~n443 & ~n458;
  assign n461 = ~n459 & n460;
  assign n462 = ~n444 & ~n461;
  assign n463 = n386 & n443;
  assign n464 = n413 & ~n447;
  assign n465 = ~n413 & n447;
  assign n466 = ~n464 & ~n465;
  assign n467 = ~n443 & n466;
  assign n468 = ~n463 & ~n467;
  assign n469 = pi04 & n468;
  assign n470 = ~pi09 & n462;
  assign n471 = pi09 & ~n462;
  assign n472 = ~n470 & ~n471;
  assign n473 = ~n394 & n443;
  assign n474 = ~n414 & ~n451;
  assign n475 = n414 & n451;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n443 & n476;
  assign n478 = ~n473 & ~n477;
  assign n479 = pi06 & ~n478;
  assign n480 = ~pi06 & n478;
  assign n481 = ~n479 & ~n480;
  assign n482 = n371 & n443;
  assign n483 = ~n416 & ~n453;
  assign n484 = n416 & n453;
  assign n485 = ~n483 & ~n484;
  assign n486 = ~n443 & n485;
  assign n487 = ~n482 & ~n486;
  assign n488 = ~pi07 & ~n487;
  assign n489 = pi07 & n487;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n411 & ~n455;
  assign n492 = n411 & n455;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n443 & ~n493;
  assign n495 = ~n364 & n443;
  assign n496 = ~n494 & ~n495;
  assign n497 = pi08 & n496;
  assign n498 = ~pi08 & ~n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n378 & n443;
  assign n501 = n415 & ~n449;
  assign n502 = ~n415 & n449;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n443 & n503;
  assign n505 = ~n500 & ~n504;
  assign n506 = pi05 & n505;
  assign n507 = ~pi05 & ~n505;
  assign n508 = ~n506 & ~n507;
  assign n509 = ~pi04 & ~n468;
  assign n510 = n83 & n87;
  assign n511 = ~n509 & n510;
  assign n512 = n481 & n511;
  assign n513 = n490 & n508;
  assign n514 = n512 & n513;
  assign n515 = n499 & n514;
  assign n516 = n472 & n515;
  assign n517 = ~n469 & n516;
  assign n518 = ~n440 & ~n445;
  assign n519 = n440 & n445;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n443 & ~n520;
  assign n522 = ~n431 & n443;
  assign n523 = ~n521 & ~n522;
  assign n524 = pi03 & n523;
  assign n525 = ~pi03 & ~n523;
  assign n526 = pi00 & ~n334;
  assign n527 = n336 & n429;
  assign n528 = ~pi01 & ~n527;
  assign n529 = n526 & n528;
  assign n530 = pi01 & ~n526;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n443 & n531;
  assign n533 = ~n434 & n443;
  assign n534 = ~n532 & ~n533;
  assign n535 = pi02 & ~n534;
  assign n536 = pi00 & ~n443;
  assign n537 = ~pi01 & n536;
  assign n538 = ~n535 & n537;
  assign n539 = ~pi02 & n534;
  assign n540 = ~n525 & ~n539;
  assign n541 = ~n538 & n540;
  assign n542 = ~n524 & ~n541;
  assign n543 = n517 & n542;
  assign n544 = ~n479 & ~n506;
  assign n545 = ~n480 & ~n488;
  assign n546 = ~n544 & n545;
  assign n547 = ~n489 & ~n497;
  assign n548 = ~n546 & n547;
  assign n549 = ~n470 & ~n498;
  assign n550 = ~n548 & n549;
  assign n551 = ~n471 & n510;
  assign n552 = ~n516 & n551;
  assign n553 = ~n550 & n552;
  assign n554 = ~n543 & ~n553;
  assign n555 = ~n535 & ~n539;
  assign n556 = ~n524 & ~n525;
  assign n557 = n84 & n555;
  assign n558 = n556 & n557;
  assign n559 = n517 & n558;
  assign n560 = n554 & ~n559;
  assign n561 = ~n462 & n560;
  assign n562 = ~n84 & ~n537;
  assign n563 = ~n539 & n562;
  assign n564 = ~n535 & ~n563;
  assign n565 = ~n525 & ~n564;
  assign n566 = ~n524 & ~n565;
  assign n567 = ~n509 & ~n566;
  assign n568 = ~n469 & ~n567;
  assign n569 = ~n506 & n568;
  assign n570 = ~n507 & ~n569;
  assign n571 = ~n480 & n570;
  assign n572 = ~n479 & ~n571;
  assign n573 = ~n489 & n572;
  assign n574 = ~n488 & ~n573;
  assign n575 = ~n497 & ~n574;
  assign n576 = ~n498 & ~n575;
  assign n577 = ~n472 & ~n576;
  assign n578 = n472 & n576;
  assign n579 = ~n560 & ~n577;
  assign n580 = ~n578 & n579;
  assign n581 = ~n561 & ~n580;
  assign n582 = ~n469 & ~n509;
  assign n583 = ~n566 & ~n582;
  assign n584 = n566 & n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n560 & ~n585;
  assign n587 = n468 & n560;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~pi05 & n588;
  assign n590 = pi10 & ~n581;
  assign n591 = ~pi10 & n581;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n499 & ~n574;
  assign n594 = n499 & n574;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n560 & ~n595;
  assign n597 = ~n496 & n560;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~pi09 & ~n598;
  assign n600 = pi09 & n598;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n478 & n560;
  assign n603 = ~n481 & ~n570;
  assign n604 = n481 & n570;
  assign n605 = ~n560 & ~n603;
  assign n606 = ~n604 & n605;
  assign n607 = ~n602 & ~n606;
  assign n608 = ~pi07 & n607;
  assign n609 = pi07 & ~n607;
  assign n610 = ~n608 & ~n609;
  assign n611 = n487 & n560;
  assign n612 = n490 & ~n572;
  assign n613 = ~n490 & n572;
  assign n614 = ~n560 & ~n612;
  assign n615 = ~n613 & n614;
  assign n616 = ~n611 & ~n615;
  assign n617 = pi08 & ~n616;
  assign n618 = ~pi08 & n616;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~pi11 & n83;
  assign n621 = n505 & n560;
  assign n622 = n508 & ~n568;
  assign n623 = ~n508 & n568;
  assign n624 = ~n622 & ~n623;
  assign n625 = ~n560 & n624;
  assign n626 = ~n621 & ~n625;
  assign n627 = pi06 & ~n626;
  assign n628 = ~pi06 & n626;
  assign n629 = ~n627 & ~n628;
  assign n630 = n620 & n629;
  assign n631 = n610 & n630;
  assign n632 = n619 & n631;
  assign n633 = n601 & n632;
  assign n634 = n592 & n633;
  assign n635 = ~n589 & n634;
  assign n636 = ~n609 & ~n627;
  assign n637 = ~n608 & ~n636;
  assign n638 = ~n618 & n637;
  assign n639 = ~n617 & ~n638;
  assign n640 = ~n600 & n639;
  assign n641 = ~n599 & ~n640;
  assign n642 = ~n591 & n641;
  assign n643 = ~n590 & n620;
  assign n644 = ~n642 & n643;
  assign n645 = ~n635 & n644;
  assign n646 = pi05 & ~n588;
  assign n647 = ~n589 & ~n646;
  assign n648 = n634 & n647;
  assign n649 = n523 & n560;
  assign n650 = n556 & ~n564;
  assign n651 = ~n556 & n564;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~n560 & n652;
  assign n654 = ~n649 & ~n653;
  assign n655 = pi04 & ~n654;
  assign n656 = ~pi04 & n654;
  assign n657 = ~n534 & n560;
  assign n658 = ~n555 & ~n562;
  assign n659 = n555 & n562;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n560 & n660;
  assign n662 = ~n657 & ~n661;
  assign n663 = pi03 & ~n662;
  assign n664 = pi00 & n439;
  assign n665 = n314 & ~n664;
  assign n666 = ~n314 & n664;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n560 & ~n667;
  assign n669 = n536 & n560;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~pi02 & ~n670;
  assign n672 = pi02 & n670;
  assign n673 = pi00 & ~n560;
  assign n674 = ~pi01 & n673;
  assign n675 = ~n672 & n674;
  assign n676 = ~pi03 & n662;
  assign n677 = ~n671 & ~n676;
  assign n678 = ~n675 & n677;
  assign n679 = ~n663 & ~n678;
  assign n680 = ~n656 & ~n679;
  assign n681 = ~n655 & ~n680;
  assign n682 = n648 & n681;
  assign n683 = ~n645 & ~n682;
  assign n684 = ~n671 & ~n672;
  assign n685 = ~n655 & ~n656;
  assign n686 = ~n663 & ~n676;
  assign n687 = n84 & n684;
  assign n688 = n685 & n686;
  assign n689 = n687 & n688;
  assign n690 = n648 & n689;
  assign n691 = n683 & ~n690;
  assign n692 = ~n581 & n691;
  assign n693 = ~n84 & ~n674;
  assign n694 = ~n672 & ~n693;
  assign n695 = ~n671 & ~n694;
  assign n696 = ~n663 & ~n695;
  assign n697 = ~n676 & ~n696;
  assign n698 = ~n655 & ~n697;
  assign n699 = ~n656 & ~n698;
  assign n700 = ~n646 & ~n699;
  assign n701 = ~n589 & ~n700;
  assign n702 = ~n627 & ~n701;
  assign n703 = ~n628 & ~n702;
  assign n704 = ~n608 & n703;
  assign n705 = ~n609 & ~n704;
  assign n706 = ~n618 & ~n705;
  assign n707 = ~n617 & ~n706;
  assign n708 = ~n599 & ~n707;
  assign n709 = ~n600 & ~n708;
  assign n710 = n592 & ~n709;
  assign n711 = ~n592 & n709;
  assign n712 = ~n691 & ~n710;
  assign n713 = ~n711 & n712;
  assign n714 = ~n692 & ~n713;
  assign n715 = ~pi11 & n714;
  assign n716 = n598 & n691;
  assign n717 = n601 & ~n707;
  assign n718 = ~n601 & n707;
  assign n719 = ~n691 & ~n717;
  assign n720 = ~n718 & n719;
  assign n721 = ~n716 & ~n720;
  assign n722 = pi10 & ~n721;
  assign n723 = pi11 & ~n714;
  assign n724 = ~pi10 & n721;
  assign n725 = ~n616 & n691;
  assign n726 = n619 & ~n705;
  assign n727 = ~n619 & n705;
  assign n728 = ~n691 & ~n726;
  assign n729 = ~n727 & n728;
  assign n730 = ~n725 & ~n729;
  assign n731 = ~pi09 & n730;
  assign n732 = ~n607 & n691;
  assign n733 = ~n610 & ~n703;
  assign n734 = n610 & n703;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~n691 & n735;
  assign n737 = ~n732 & ~n736;
  assign n738 = pi08 & ~n737;
  assign n739 = ~pi08 & n737;
  assign n740 = ~n738 & ~n739;
  assign n741 = n588 & n691;
  assign n742 = n647 & ~n699;
  assign n743 = ~n647 & n699;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n691 & n744;
  assign n746 = ~n741 & ~n745;
  assign n747 = ~pi06 & ~n746;
  assign n748 = ~n626 & n691;
  assign n749 = ~n629 & ~n701;
  assign n750 = n629 & n701;
  assign n751 = ~n749 & ~n750;
  assign n752 = ~n691 & n751;
  assign n753 = ~n748 & ~n752;
  assign n754 = pi07 & ~n753;
  assign n755 = ~pi07 & n753;
  assign n756 = ~n754 & ~n755;
  assign n757 = n83 & ~n747;
  assign n758 = n740 & n757;
  assign n759 = n756 & n758;
  assign n760 = pi09 & ~n730;
  assign n761 = ~n739 & n754;
  assign n762 = ~n738 & ~n760;
  assign n763 = ~n761 & n762;
  assign n764 = ~n759 & n763;
  assign n765 = ~n724 & ~n731;
  assign n766 = ~n764 & n765;
  assign n767 = ~n722 & ~n723;
  assign n768 = ~n766 & n767;
  assign n769 = ~n715 & ~n768;
  assign n770 = n83 & ~n769;
  assign n771 = pi06 & n746;
  assign n772 = ~n731 & ~n760;
  assign n773 = ~n715 & ~n723;
  assign n774 = ~n722 & ~n724;
  assign n775 = ~n771 & n772;
  assign n776 = n759 & n775;
  assign n777 = n774 & n776;
  assign n778 = n773 & n777;
  assign n779 = n654 & n691;
  assign n780 = n685 & ~n697;
  assign n781 = ~n685 & n697;
  assign n782 = ~n780 & ~n781;
  assign n783 = ~n691 & n782;
  assign n784 = ~n779 & ~n783;
  assign n785 = pi05 & n784;
  assign n786 = ~pi05 & ~n784;
  assign n787 = n662 & n691;
  assign n788 = n686 & ~n695;
  assign n789 = ~n686 & n695;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n691 & n790;
  assign n792 = ~n787 & ~n791;
  assign n793 = pi04 & n792;
  assign n794 = ~n684 & ~n693;
  assign n795 = n684 & n693;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~n691 & ~n796;
  assign n798 = ~n670 & n691;
  assign n799 = ~n797 & ~n798;
  assign n800 = pi03 & n799;
  assign n801 = n314 & n554;
  assign n802 = pi01 & ~n554;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n691 & n803;
  assign n805 = ~n673 & n691;
  assign n806 = ~n804 & ~n805;
  assign n807 = pi02 & ~n806;
  assign n808 = ~n800 & ~n807;
  assign n809 = ~pi03 & ~n799;
  assign n810 = ~pi04 & ~n792;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n808 & n811;
  assign n813 = ~n793 & ~n812;
  assign n814 = ~n786 & ~n813;
  assign n815 = ~n785 & ~n814;
  assign n816 = n778 & n815;
  assign n817 = ~n770 & ~n816;
  assign n818 = ~n785 & ~n786;
  assign n819 = ~n793 & ~n810;
  assign n820 = ~n800 & ~n809;
  assign n821 = ~pi02 & n806;
  assign n822 = ~n807 & ~n821;
  assign n823 = n818 & n819;
  assign n824 = n820 & n822;
  assign n825 = n823 & n824;
  assign n826 = n778 & n825;
  assign n827 = ~n817 & ~n826;
  assign n828 = pi00 & n691;
  assign n829 = ~pi01 & ~n828;
  assign n830 = n826 & n829;
  assign n831 = ~n827 & ~n830;
  assign n832 = ~n747 & ~n771;
  assign n833 = ~n821 & ~n829;
  assign n834 = ~n807 & ~n833;
  assign n835 = ~n800 & n834;
  assign n836 = ~n809 & ~n835;
  assign n837 = ~n810 & n836;
  assign n838 = ~n793 & ~n837;
  assign n839 = ~n785 & n838;
  assign n840 = ~n786 & ~n839;
  assign n841 = ~n832 & n840;
  assign n842 = ~n771 & ~n840;
  assign n843 = ~n747 & n842;
  assign n844 = ~n841 & ~n843;
  assign n845 = ~n831 & ~n844;
  assign n846 = n746 & n831;
  assign n847 = ~n845 & ~n846;
  assign n848 = ~n714 & n831;
  assign n849 = ~n747 & ~n842;
  assign n850 = ~n754 & ~n849;
  assign n851 = ~n755 & ~n850;
  assign n852 = ~n739 & n851;
  assign n853 = ~n738 & ~n852;
  assign n854 = ~n731 & ~n853;
  assign n855 = ~n760 & ~n854;
  assign n856 = ~n724 & ~n855;
  assign n857 = ~n722 & ~n856;
  assign n858 = n773 & ~n857;
  assign n859 = ~n773 & n857;
  assign n860 = ~n831 & ~n858;
  assign n861 = ~n859 & n860;
  assign n862 = ~n848 & ~n861;
  assign n863 = ~pi12 & n862;
  assign n864 = pi12 & ~n862;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~n730 & n831;
  assign n867 = n772 & ~n853;
  assign n868 = ~n772 & n853;
  assign n869 = ~n831 & ~n867;
  assign n870 = ~n868 & n869;
  assign n871 = ~n866 & ~n870;
  assign n872 = ~pi10 & n871;
  assign n873 = pi10 & ~n871;
  assign n874 = ~n872 & ~n873;
  assign n875 = pi07 & ~n847;
  assign n876 = ~n721 & n831;
  assign n877 = n774 & ~n855;
  assign n878 = ~n774 & n855;
  assign n879 = ~n831 & ~n877;
  assign n880 = ~n878 & n879;
  assign n881 = ~n876 & ~n880;
  assign n882 = pi11 & ~n881;
  assign n883 = ~pi11 & n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n737 & n831;
  assign n886 = ~n740 & ~n851;
  assign n887 = n740 & n851;
  assign n888 = ~n831 & ~n886;
  assign n889 = ~n887 & n888;
  assign n890 = ~n885 & ~n889;
  assign n891 = pi09 & ~n890;
  assign n892 = ~pi09 & n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~pi07 & n847;
  assign n895 = n753 & n831;
  assign n896 = n756 & ~n849;
  assign n897 = ~n756 & n849;
  assign n898 = ~n896 & ~n897;
  assign n899 = ~n831 & n898;
  assign n900 = ~n895 & ~n899;
  assign n901 = pi08 & n900;
  assign n902 = ~pi08 & ~n900;
  assign n903 = ~n901 & ~n902;
  assign n904 = n82 & ~n894;
  assign n905 = n903 & n904;
  assign n906 = ~n875 & n905;
  assign n907 = n893 & n906;
  assign n908 = n874 & n907;
  assign n909 = n884 & n908;
  assign n910 = n865 & n909;
  assign n911 = ~n818 & ~n838;
  assign n912 = n818 & n838;
  assign n913 = ~n911 & ~n912;
  assign n914 = ~n831 & ~n913;
  assign n915 = n784 & n831;
  assign n916 = ~n914 & ~n915;
  assign n917 = ~pi06 & n916;
  assign n918 = pi06 & ~n916;
  assign n919 = ~n819 & ~n836;
  assign n920 = n819 & n836;
  assign n921 = ~n919 & ~n920;
  assign n922 = ~n831 & ~n921;
  assign n923 = ~n792 & n831;
  assign n924 = ~n922 & ~n923;
  assign n925 = pi05 & n924;
  assign n926 = n799 & n831;
  assign n927 = n820 & ~n834;
  assign n928 = ~n820 & n834;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n831 & n929;
  assign n931 = ~n926 & ~n930;
  assign n932 = ~pi04 & n931;
  assign n933 = ~pi05 & ~n924;
  assign n934 = n806 & n831;
  assign n935 = ~n822 & ~n829;
  assign n936 = n822 & n829;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n831 & n937;
  assign n939 = ~n934 & ~n938;
  assign n940 = pi03 & n939;
  assign n941 = pi04 & ~n931;
  assign n942 = ~n940 & ~n941;
  assign n943 = ~n932 & ~n933;
  assign n944 = ~n942 & n943;
  assign n945 = ~n918 & ~n925;
  assign n946 = ~n944 & n945;
  assign n947 = ~n917 & ~n946;
  assign n948 = n910 & ~n947;
  assign n949 = ~n891 & ~n901;
  assign n950 = ~n905 & n949;
  assign n951 = ~n872 & ~n892;
  assign n952 = ~n950 & n951;
  assign n953 = ~n873 & ~n882;
  assign n954 = ~n952 & n953;
  assign n955 = ~n863 & ~n883;
  assign n956 = ~n954 & n955;
  assign n957 = n82 & ~n864;
  assign n958 = ~n956 & n957;
  assign n959 = ~n948 & ~n958;
  assign n960 = pi00 & ~n691;
  assign n961 = n831 & ~n960;
  assign n962 = n314 & n683;
  assign n963 = pi01 & ~n683;
  assign n964 = ~n962 & ~n963;
  assign n965 = ~n831 & n964;
  assign n966 = ~n961 & ~n965;
  assign n967 = pi02 & ~n966;
  assign n968 = ~pi02 & n966;
  assign n969 = pi00 & ~n831;
  assign n970 = ~pi01 & n969;
  assign n971 = ~n968 & ~n970;
  assign n972 = ~n967 & ~n971;
  assign n973 = ~n932 & ~n941;
  assign n974 = ~n917 & ~n918;
  assign n975 = ~n925 & ~n933;
  assign n976 = ~pi03 & ~n939;
  assign n977 = ~n940 & ~n976;
  assign n978 = n973 & n974;
  assign n979 = n975 & n977;
  assign n980 = n978 & n979;
  assign n981 = n910 & n980;
  assign n982 = ~n972 & n981;
  assign n983 = ~n959 & ~n982;
  assign n984 = ~n967 & ~n968;
  assign n985 = n84 & n984;
  assign n986 = n981 & n985;
  assign n987 = ~n983 & ~n986;
  assign n988 = ~n847 & n987;
  assign n989 = ~n84 & ~n970;
  assign n990 = ~n967 & ~n989;
  assign n991 = ~n968 & ~n990;
  assign n992 = ~n940 & ~n991;
  assign n993 = ~n976 & ~n992;
  assign n994 = ~n932 & n993;
  assign n995 = ~n941 & ~n994;
  assign n996 = ~n933 & ~n995;
  assign n997 = ~n925 & ~n996;
  assign n998 = ~n917 & ~n997;
  assign n999 = ~n918 & ~n998;
  assign n1000 = ~n875 & ~n894;
  assign n1001 = n999 & ~n1000;
  assign n1002 = ~n999 & n1000;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~n987 & n1003;
  assign n1005 = ~n988 & ~n1004;
  assign n1006 = ~n862 & n987;
  assign n1007 = ~n894 & ~n999;
  assign n1008 = ~n875 & ~n1007;
  assign n1009 = ~n902 & ~n1008;
  assign n1010 = ~n901 & ~n1009;
  assign n1011 = ~n891 & n1010;
  assign n1012 = ~n892 & ~n1011;
  assign n1013 = ~n872 & n1012;
  assign n1014 = ~n873 & ~n1013;
  assign n1015 = ~n883 & ~n1014;
  assign n1016 = ~n882 & ~n1015;
  assign n1017 = n865 & ~n1016;
  assign n1018 = ~n865 & n1016;
  assign n1019 = ~n987 & ~n1017;
  assign n1020 = ~n1018 & n1019;
  assign n1021 = ~n1006 & ~n1020;
  assign n1022 = pi13 & ~n1021;
  assign n1023 = ~pi13 & n1021;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n881 & n987;
  assign n1026 = n884 & ~n1014;
  assign n1027 = ~n884 & n1014;
  assign n1028 = ~n987 & ~n1026;
  assign n1029 = ~n1027 & n1028;
  assign n1030 = ~n1025 & ~n1029;
  assign n1031 = pi12 & ~n1030;
  assign n1032 = ~pi12 & n1030;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = n890 & n987;
  assign n1035 = ~n893 & ~n1010;
  assign n1036 = n893 & n1010;
  assign n1037 = ~n987 & ~n1035;
  assign n1038 = ~n1036 & n1037;
  assign n1039 = ~n1034 & ~n1038;
  assign n1040 = pi10 & n1039;
  assign n1041 = ~pi10 & ~n1039;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = pi08 & ~n1005;
  assign n1044 = ~pi08 & n1005;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~n903 & ~n1008;
  assign n1047 = n903 & n1008;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n987 & ~n1048;
  assign n1050 = n900 & n987;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = pi09 & ~n1051;
  assign n1053 = ~pi09 & n1051;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = n81 & n1054;
  assign n1056 = ~n871 & n987;
  assign n1057 = ~n874 & ~n1012;
  assign n1058 = n874 & n1012;
  assign n1059 = ~n987 & ~n1057;
  assign n1060 = ~n1058 & n1059;
  assign n1061 = ~n1056 & ~n1060;
  assign n1062 = pi11 & ~n1061;
  assign n1063 = ~pi11 & n1061;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n1045 & n1055;
  assign n1066 = n1042 & n1065;
  assign n1067 = n1064 & n1066;
  assign n1068 = n1033 & n1067;
  assign n1069 = n1024 & n1068;
  assign n1070 = n931 & n987;
  assign n1071 = n973 & ~n993;
  assign n1072 = ~n973 & n993;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = ~n987 & n1073;
  assign n1075 = ~n1070 & ~n1074;
  assign n1076 = pi05 & n1075;
  assign n1077 = ~pi05 & ~n1075;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~n916 & n987;
  assign n1080 = n974 & ~n997;
  assign n1081 = ~n974 & n997;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = ~n987 & n1082;
  assign n1084 = ~n1079 & ~n1083;
  assign n1085 = pi07 & ~n1084;
  assign n1086 = ~pi07 & n1084;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = n924 & n987;
  assign n1089 = n975 & ~n995;
  assign n1090 = ~n975 & n995;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n987 & n1091;
  assign n1093 = ~n1088 & ~n1092;
  assign n1094 = pi06 & ~n1093;
  assign n1095 = ~pi06 & n1093;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n939 & n987;
  assign n1098 = n977 & ~n991;
  assign n1099 = ~n977 & n991;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~n987 & n1100;
  assign n1102 = ~n1097 & ~n1101;
  assign n1103 = pi04 & n1102;
  assign n1104 = ~pi04 & ~n1102;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = n1078 & n1087;
  assign n1107 = n1096 & n1105;
  assign n1108 = n1106 & n1107;
  assign n1109 = n1069 & n1108;
  assign n1110 = ~n966 & n987;
  assign n1111 = ~n984 & ~n989;
  assign n1112 = n984 & n989;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n987 & n1113;
  assign n1115 = ~n1110 & ~n1114;
  assign n1116 = pi03 & ~n1115;
  assign n1117 = pi00 & ~n827;
  assign n1118 = n826 & n960;
  assign n1119 = ~pi01 & ~n1118;
  assign n1120 = n1117 & n1119;
  assign n1121 = pi01 & ~n1117;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = ~n987 & n1122;
  assign n1124 = ~n969 & n987;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~pi02 & n1125;
  assign n1127 = pi00 & ~n987;
  assign n1128 = ~pi01 & n1127;
  assign n1129 = pi02 & ~n1125;
  assign n1130 = n1128 & ~n1129;
  assign n1131 = ~pi03 & n1115;
  assign n1132 = ~n1126 & ~n1131;
  assign n1133 = ~n1130 & n1132;
  assign n1134 = ~n1116 & ~n1133;
  assign n1135 = n1109 & ~n1134;
  assign n1136 = ~n1077 & n1103;
  assign n1137 = ~n1076 & ~n1094;
  assign n1138 = ~n1136 & n1137;
  assign n1139 = ~n1086 & ~n1095;
  assign n1140 = ~n1138 & n1139;
  assign n1141 = ~n1085 & ~n1140;
  assign n1142 = n1069 & n1141;
  assign n1143 = ~n1044 & n1055;
  assign n1144 = ~n1040 & ~n1052;
  assign n1145 = ~n1143 & n1144;
  assign n1146 = ~n1041 & ~n1063;
  assign n1147 = ~n1145 & n1146;
  assign n1148 = ~n1031 & ~n1062;
  assign n1149 = ~n1147 & n1148;
  assign n1150 = ~n1023 & ~n1032;
  assign n1151 = ~n1149 & n1150;
  assign n1152 = n81 & ~n1022;
  assign n1153 = ~n1151 & n1152;
  assign n1154 = ~n1142 & ~n1153;
  assign n1155 = ~n1135 & ~n1154;
  assign n1156 = ~n1116 & ~n1131;
  assign n1157 = ~n1126 & ~n1129;
  assign n1158 = n84 & n1156;
  assign n1159 = n1157 & n1158;
  assign n1160 = n1109 & n1159;
  assign n1161 = ~n1155 & ~n1160;
  assign n1162 = n1005 & n1161;
  assign n1163 = ~n84 & ~n1128;
  assign n1164 = ~n1126 & n1163;
  assign n1165 = ~n1129 & ~n1164;
  assign n1166 = ~n1131 & ~n1165;
  assign n1167 = ~n1116 & ~n1166;
  assign n1168 = ~n1103 & n1167;
  assign n1169 = ~n1104 & ~n1168;
  assign n1170 = ~n1076 & ~n1169;
  assign n1171 = ~n1077 & ~n1170;
  assign n1172 = ~n1095 & n1171;
  assign n1173 = ~n1094 & ~n1172;
  assign n1174 = ~n1086 & ~n1173;
  assign n1175 = ~n1085 & ~n1174;
  assign n1176 = ~n1045 & ~n1175;
  assign n1177 = n1045 & n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1161 & n1178;
  assign n1180 = ~n1162 & ~n1179;
  assign n1181 = ~n1115 & n1161;
  assign n1182 = n1156 & ~n1165;
  assign n1183 = ~n1156 & n1165;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n1161 & n1184;
  assign n1186 = ~n1181 & ~n1185;
  assign n1187 = pi04 & ~n1186;
  assign n1188 = ~pi04 & n1186;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1125 & n1161;
  assign n1191 = ~n1157 & ~n1163;
  assign n1192 = n1157 & n1163;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1161 & n1193;
  assign n1195 = ~n1190 & ~n1194;
  assign n1196 = pi03 & ~n1195;
  assign n1197 = ~pi03 & n1195;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = n1093 & n1161;
  assign n1200 = n1096 & ~n1171;
  assign n1201 = ~n1096 & n1171;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1161 & n1202;
  assign n1204 = ~n1199 & ~n1203;
  assign n1205 = pi07 & n1204;
  assign n1206 = ~pi07 & ~n1204;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~n1075 & n1161;
  assign n1209 = n1078 & ~n1169;
  assign n1210 = ~n1078 & n1169;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1161 & n1211;
  assign n1213 = ~n1208 & ~n1212;
  assign n1214 = pi06 & n1213;
  assign n1215 = ~pi06 & ~n1213;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1084 & n1161;
  assign n1218 = n1087 & ~n1173;
  assign n1219 = ~n1087 & n1173;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = ~n1161 & n1220;
  assign n1222 = ~n1217 & ~n1221;
  assign n1223 = pi08 & ~n1222;
  assign n1224 = ~pi08 & n1222;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = ~pi09 & ~n1180;
  assign n1227 = pi09 & n1180;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n1021 & n1161;
  assign n1230 = ~n1044 & ~n1175;
  assign n1231 = ~n1043 & ~n1230;
  assign n1232 = ~n1053 & ~n1231;
  assign n1233 = ~n1052 & ~n1232;
  assign n1234 = ~n1040 & n1233;
  assign n1235 = ~n1041 & ~n1234;
  assign n1236 = ~n1063 & n1235;
  assign n1237 = ~n1062 & ~n1236;
  assign n1238 = ~n1032 & ~n1237;
  assign n1239 = ~n1031 & ~n1238;
  assign n1240 = n1024 & ~n1239;
  assign n1241 = ~n1024 & n1239;
  assign n1242 = ~n1161 & ~n1240;
  assign n1243 = ~n1241 & n1242;
  assign n1244 = ~n1229 & ~n1243;
  assign n1245 = pi14 & ~n1244;
  assign n1246 = ~pi14 & n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n1061 & n1161;
  assign n1249 = ~n1064 & ~n1235;
  assign n1250 = n1064 & n1235;
  assign n1251 = ~n1161 & ~n1249;
  assign n1252 = ~n1250 & n1251;
  assign n1253 = ~n1248 & ~n1252;
  assign n1254 = pi12 & ~n1253;
  assign n1255 = ~pi12 & n1253;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n1030 & n1161;
  assign n1258 = n1033 & ~n1237;
  assign n1259 = ~n1033 & n1237;
  assign n1260 = ~n1161 & ~n1258;
  assign n1261 = ~n1259 & n1260;
  assign n1262 = ~n1257 & ~n1261;
  assign n1263 = pi13 & ~n1262;
  assign n1264 = ~pi13 & n1262;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = n1039 & n1161;
  assign n1267 = n1042 & ~n1233;
  assign n1268 = ~n1042 & n1233;
  assign n1269 = ~n1161 & ~n1267;
  assign n1270 = ~n1268 & n1269;
  assign n1271 = ~n1266 & ~n1270;
  assign n1272 = pi11 & ~n1271;
  assign n1273 = ~pi11 & n1271;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1051 & n1161;
  assign n1276 = n1054 & ~n1231;
  assign n1277 = ~n1054 & n1231;
  assign n1278 = ~n1161 & ~n1276;
  assign n1279 = ~n1277 & n1278;
  assign n1280 = ~n1275 & ~n1279;
  assign n1281 = pi10 & ~n1280;
  assign n1282 = ~pi10 & n1280;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = n80 & n1283;
  assign n1285 = n1274 & n1284;
  assign n1286 = n1256 & n1285;
  assign n1287 = n1265 & n1286;
  assign n1288 = n1247 & n1287;
  assign n1289 = n1228 & n1288;
  assign n1290 = n1102 & n1161;
  assign n1291 = n1105 & ~n1167;
  assign n1292 = ~n1105 & n1167;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1161 & n1293;
  assign n1295 = ~n1290 & ~n1294;
  assign n1296 = pi05 & ~n1295;
  assign n1297 = ~pi05 & n1295;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = n1207 & n1216;
  assign n1300 = n1225 & n1298;
  assign n1301 = n1299 & n1300;
  assign n1302 = n1289 & n1301;
  assign n1303 = n1189 & n1198;
  assign n1304 = n1302 & n1303;
  assign n1305 = pi01 & n983;
  assign n1306 = n314 & ~n983;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1161 & n1307;
  assign n1309 = ~n1127 & n1161;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = pi02 & ~n1310;
  assign n1312 = ~pi02 & n1310;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = pi00 & ~n1161;
  assign n1315 = ~pi01 & n1314;
  assign n1316 = n1313 & ~n1315;
  assign n1317 = n1304 & n1316;
  assign n1318 = ~n1226 & n1288;
  assign n1319 = ~n1272 & ~n1281;
  assign n1320 = ~n1273 & ~n1319;
  assign n1321 = ~n1255 & n1320;
  assign n1322 = ~n1254 & ~n1321;
  assign n1323 = ~n1263 & n1322;
  assign n1324 = ~n1264 & ~n1323;
  assign n1325 = ~n1246 & n1324;
  assign n1326 = n80 & ~n1245;
  assign n1327 = ~n1325 & n1326;
  assign n1328 = ~n1318 & n1327;
  assign n1329 = ~n1215 & n1296;
  assign n1330 = ~n1205 & ~n1214;
  assign n1331 = ~n1329 & n1330;
  assign n1332 = ~n1206 & ~n1331;
  assign n1333 = ~n1223 & ~n1332;
  assign n1334 = ~n1224 & ~n1333;
  assign n1335 = n1289 & ~n1334;
  assign n1336 = ~n1328 & ~n1335;
  assign n1337 = ~n1302 & ~n1336;
  assign n1338 = ~n1197 & n1311;
  assign n1339 = ~n1187 & ~n1196;
  assign n1340 = ~n1338 & n1339;
  assign n1341 = ~n1188 & ~n1340;
  assign n1342 = n1302 & ~n1341;
  assign n1343 = ~n1337 & ~n1342;
  assign n1344 = ~n1317 & ~n1343;
  assign n1345 = n84 & n1313;
  assign n1346 = n1304 & n1345;
  assign n1347 = ~n1344 & ~n1346;
  assign n1348 = n1180 & n1347;
  assign n1349 = ~n84 & ~n1315;
  assign n1350 = ~n1311 & ~n1349;
  assign n1351 = ~n1312 & ~n1350;
  assign n1352 = ~n1197 & n1351;
  assign n1353 = ~n1196 & ~n1352;
  assign n1354 = ~n1188 & ~n1353;
  assign n1355 = ~n1187 & ~n1354;
  assign n1356 = ~n1297 & ~n1355;
  assign n1357 = ~n1296 & ~n1356;
  assign n1358 = ~n1215 & ~n1357;
  assign n1359 = ~n1214 & ~n1358;
  assign n1360 = ~n1206 & ~n1359;
  assign n1361 = ~n1205 & ~n1360;
  assign n1362 = ~n1224 & ~n1361;
  assign n1363 = ~n1223 & ~n1362;
  assign n1364 = n1228 & ~n1363;
  assign n1365 = ~n1228 & n1363;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1347 & n1366;
  assign n1368 = ~n1348 & ~n1367;
  assign n1369 = pi10 & ~n1368;
  assign n1370 = ~n1262 & n1347;
  assign n1371 = ~n1226 & ~n1363;
  assign n1372 = ~n1227 & ~n1371;
  assign n1373 = ~n1282 & ~n1372;
  assign n1374 = ~n1281 & ~n1373;
  assign n1375 = ~n1272 & n1374;
  assign n1376 = ~n1273 & ~n1375;
  assign n1377 = ~n1255 & n1376;
  assign n1378 = ~n1254 & ~n1377;
  assign n1379 = n1265 & ~n1378;
  assign n1380 = ~n1265 & n1378;
  assign n1381 = ~n1347 & ~n1379;
  assign n1382 = ~n1380 & n1381;
  assign n1383 = ~n1370 & ~n1382;
  assign n1384 = pi14 & ~n1383;
  assign n1385 = ~pi14 & n1383;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n1271 & n1347;
  assign n1388 = n1274 & ~n1374;
  assign n1389 = ~n1274 & n1374;
  assign n1390 = ~n1347 & ~n1388;
  assign n1391 = ~n1389 & n1390;
  assign n1392 = ~n1387 & ~n1391;
  assign n1393 = pi12 & ~n1392;
  assign n1394 = ~pi12 & n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = ~n1244 & n1347;
  assign n1397 = ~n1264 & ~n1378;
  assign n1398 = ~n1263 & ~n1397;
  assign n1399 = n1247 & ~n1398;
  assign n1400 = ~n1247 & n1398;
  assign n1401 = ~n1347 & ~n1399;
  assign n1402 = ~n1400 & n1401;
  assign n1403 = ~n1396 & ~n1402;
  assign n1404 = pi15 & ~n1403;
  assign n1405 = ~pi15 & n1403;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = ~n1253 & n1347;
  assign n1408 = ~n1256 & ~n1376;
  assign n1409 = n1256 & n1376;
  assign n1410 = ~n1347 & ~n1408;
  assign n1411 = ~n1409 & n1410;
  assign n1412 = ~n1407 & ~n1411;
  assign n1413 = pi13 & ~n1412;
  assign n1414 = ~pi13 & n1412;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~pi18 & n76;
  assign n1417 = ~pi17 & n1416;
  assign n1418 = ~pi16 & n1417;
  assign n1419 = n1280 & n1347;
  assign n1420 = ~n1283 & ~n1372;
  assign n1421 = n1283 & n1372;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1347 & n1422;
  assign n1424 = ~n1419 & ~n1423;
  assign n1425 = pi11 & n1424;
  assign n1426 = ~pi11 & ~n1424;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~pi10 & n1368;
  assign n1429 = n1418 & ~n1428;
  assign n1430 = n1427 & n1429;
  assign n1431 = n1395 & n1430;
  assign n1432 = n1415 & n1431;
  assign n1433 = n1386 & n1432;
  assign n1434 = n1406 & n1433;
  assign n1435 = ~n1369 & n1434;
  assign n1436 = n1204 & n1347;
  assign n1437 = n1207 & ~n1359;
  assign n1438 = ~n1207 & n1359;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~n1347 & n1439;
  assign n1441 = ~n1436 & ~n1440;
  assign n1442 = ~pi08 & n1441;
  assign n1443 = pi08 & ~n1441;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = n1213 & n1347;
  assign n1446 = n1216 & ~n1357;
  assign n1447 = ~n1216 & n1357;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1347 & n1448;
  assign n1450 = ~n1445 & ~n1449;
  assign n1451 = pi07 & ~n1450;
  assign n1452 = ~pi07 & n1450;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = ~n1222 & n1347;
  assign n1455 = n1225 & ~n1361;
  assign n1456 = ~n1225 & n1361;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n1347 & n1457;
  assign n1459 = ~n1454 & ~n1458;
  assign n1460 = pi09 & ~n1459;
  assign n1461 = ~pi09 & n1459;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = ~n1295 & n1347;
  assign n1464 = n1298 & ~n1355;
  assign n1465 = ~n1298 & n1355;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = ~n1347 & n1466;
  assign n1468 = ~n1463 & ~n1467;
  assign n1469 = pi06 & ~n1468;
  assign n1470 = ~pi06 & n1468;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = n1444 & n1453;
  assign n1473 = n1462 & n1471;
  assign n1474 = n1472 & n1473;
  assign n1475 = n1435 & n1474;
  assign n1476 = ~n1393 & ~n1425;
  assign n1477 = ~n1394 & ~n1476;
  assign n1478 = ~n1414 & n1477;
  assign n1479 = ~n1413 & ~n1478;
  assign n1480 = ~n1384 & n1479;
  assign n1481 = ~n1385 & ~n1480;
  assign n1482 = ~n1405 & n1481;
  assign n1483 = ~n1404 & n1418;
  assign n1484 = ~n1482 & n1483;
  assign n1485 = ~n1434 & n1484;
  assign n1486 = ~n1452 & n1469;
  assign n1487 = ~n1443 & ~n1451;
  assign n1488 = ~n1486 & n1487;
  assign n1489 = ~n1442 & ~n1461;
  assign n1490 = ~n1488 & n1489;
  assign n1491 = ~n1460 & ~n1490;
  assign n1492 = n1435 & n1491;
  assign n1493 = ~n1475 & ~n1485;
  assign n1494 = ~n1492 & n1493;
  assign n1495 = ~n1310 & n1347;
  assign n1496 = ~n1313 & ~n1349;
  assign n1497 = n1313 & n1349;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~n1347 & n1498;
  assign n1500 = ~n1495 & ~n1499;
  assign n1501 = pi03 & ~n1500;
  assign n1502 = ~pi03 & n1500;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~n1195 & n1347;
  assign n1505 = ~n1198 & ~n1351;
  assign n1506 = n1198 & n1351;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1347 & n1507;
  assign n1509 = ~n1504 & ~n1508;
  assign n1510 = ~pi04 & n1509;
  assign n1511 = pi04 & ~n1509;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = pi01 & n1155;
  assign n1514 = n314 & ~n1155;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~n1347 & n1515;
  assign n1517 = ~n1314 & n1347;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~pi02 & n1518;
  assign n1520 = ~n1186 & n1347;
  assign n1521 = n1189 & ~n1353;
  assign n1522 = ~n1189 & n1353;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1347 & n1523;
  assign n1525 = ~n1520 & ~n1524;
  assign n1526 = pi05 & ~n1525;
  assign n1527 = ~pi05 & n1525;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = n1503 & ~n1519;
  assign n1530 = n1512 & n1528;
  assign n1531 = n1529 & n1530;
  assign n1532 = ~n1501 & ~n1511;
  assign n1533 = ~n1510 & ~n1527;
  assign n1534 = ~n1532 & n1533;
  assign n1535 = ~n1526 & ~n1534;
  assign n1536 = ~n1531 & n1535;
  assign n1537 = n1475 & ~n1536;
  assign n1538 = ~n1494 & ~n1537;
  assign n1539 = pi00 & n1347;
  assign n1540 = ~pi01 & ~n1539;
  assign n1541 = pi02 & ~n1518;
  assign n1542 = n1531 & ~n1541;
  assign n1543 = n1475 & n1542;
  assign n1544 = n1540 & n1543;
  assign n1545 = ~n1538 & ~n1544;
  assign n1546 = pi00 & ~n1344;
  assign n1547 = ~pi01 & ~n1546;
  assign n1548 = pi01 & n1546;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1545 & ~n1549;
  assign n1551 = pi00 & ~n1347;
  assign n1552 = n1545 & ~n1551;
  assign n1553 = ~n1550 & ~n1552;
  assign n1554 = n1368 & n1545;
  assign n1555 = ~n1369 & ~n1428;
  assign n1556 = ~n1519 & ~n1540;
  assign n1557 = ~n1541 & ~n1556;
  assign n1558 = ~n1502 & ~n1557;
  assign n1559 = ~n1501 & ~n1558;
  assign n1560 = ~n1511 & n1559;
  assign n1561 = ~n1510 & ~n1560;
  assign n1562 = ~n1527 & n1561;
  assign n1563 = ~n1526 & ~n1562;
  assign n1564 = ~n1470 & ~n1563;
  assign n1565 = ~n1469 & ~n1564;
  assign n1566 = ~n1452 & ~n1565;
  assign n1567 = ~n1451 & ~n1566;
  assign n1568 = ~n1442 & ~n1567;
  assign n1569 = ~n1443 & ~n1568;
  assign n1570 = ~n1461 & ~n1569;
  assign n1571 = ~n1460 & ~n1570;
  assign n1572 = ~n1555 & ~n1571;
  assign n1573 = n1555 & n1571;
  assign n1574 = ~n1545 & ~n1572;
  assign n1575 = ~n1573 & n1574;
  assign n1576 = ~n1554 & ~n1575;
  assign n1577 = ~pi11 & ~n1576;
  assign n1578 = ~n1403 & n1545;
  assign n1579 = ~n1428 & ~n1571;
  assign n1580 = ~n1369 & ~n1579;
  assign n1581 = ~n1426 & ~n1580;
  assign n1582 = ~n1425 & ~n1581;
  assign n1583 = ~n1393 & n1582;
  assign n1584 = ~n1394 & ~n1583;
  assign n1585 = ~n1414 & n1584;
  assign n1586 = ~n1413 & ~n1585;
  assign n1587 = ~n1385 & ~n1586;
  assign n1588 = ~n1384 & ~n1587;
  assign n1589 = n1406 & ~n1588;
  assign n1590 = ~n1406 & n1588;
  assign n1591 = ~n1545 & ~n1589;
  assign n1592 = ~n1590 & n1591;
  assign n1593 = ~n1578 & ~n1592;
  assign n1594 = pi16 & ~n1593;
  assign n1595 = ~pi16 & n1593;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = ~n1427 & ~n1580;
  assign n1598 = n1427 & n1580;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~n1545 & ~n1599;
  assign n1601 = n1424 & n1545;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = pi12 & ~n1602;
  assign n1604 = ~pi12 & n1602;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = ~n1383 & n1545;
  assign n1607 = n1386 & ~n1586;
  assign n1608 = ~n1386 & n1586;
  assign n1609 = ~n1545 & ~n1607;
  assign n1610 = ~n1608 & n1609;
  assign n1611 = ~n1606 & ~n1610;
  assign n1612 = pi15 & ~n1611;
  assign n1613 = ~pi15 & n1611;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = ~n1392 & n1545;
  assign n1616 = n1395 & ~n1582;
  assign n1617 = ~n1395 & n1582;
  assign n1618 = ~n1545 & ~n1616;
  assign n1619 = ~n1617 & n1618;
  assign n1620 = ~n1615 & ~n1619;
  assign n1621 = pi13 & ~n1620;
  assign n1622 = ~pi13 & n1620;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = ~n1412 & n1545;
  assign n1625 = ~n1415 & ~n1584;
  assign n1626 = n1415 & n1584;
  assign n1627 = ~n1545 & ~n1625;
  assign n1628 = ~n1626 & n1627;
  assign n1629 = ~n1624 & ~n1628;
  assign n1630 = pi14 & ~n1629;
  assign n1631 = ~pi14 & n1629;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = n1417 & n1605;
  assign n1634 = n1623 & n1633;
  assign n1635 = n1632 & n1634;
  assign n1636 = n1614 & n1635;
  assign n1637 = n1596 & n1636;
  assign n1638 = ~n1577 & n1637;
  assign n1639 = ~n1603 & ~n1621;
  assign n1640 = ~n1622 & ~n1639;
  assign n1641 = ~n1631 & n1640;
  assign n1642 = ~n1630 & ~n1641;
  assign n1643 = ~n1612 & n1642;
  assign n1644 = ~n1613 & ~n1643;
  assign n1645 = ~n1595 & n1644;
  assign n1646 = n1417 & ~n1594;
  assign n1647 = ~n1645 & n1646;
  assign n1648 = ~n1638 & n1647;
  assign n1649 = pi11 & n1576;
  assign n1650 = ~n1577 & ~n1649;
  assign n1651 = n1637 & n1650;
  assign n1652 = ~n1459 & n1545;
  assign n1653 = n1462 & ~n1569;
  assign n1654 = ~n1462 & n1569;
  assign n1655 = ~n1545 & ~n1653;
  assign n1656 = ~n1654 & n1655;
  assign n1657 = ~n1652 & ~n1656;
  assign n1658 = pi10 & ~n1657;
  assign n1659 = ~pi10 & n1657;
  assign n1660 = ~n1441 & n1545;
  assign n1661 = n1444 & ~n1567;
  assign n1662 = ~n1444 & n1567;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = ~n1545 & n1663;
  assign n1665 = ~n1660 & ~n1664;
  assign n1666 = ~pi09 & n1665;
  assign n1667 = ~n1450 & n1545;
  assign n1668 = n1453 & ~n1565;
  assign n1669 = ~n1453 & n1565;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = ~n1545 & n1670;
  assign n1672 = ~n1667 & ~n1671;
  assign n1673 = ~pi08 & n1672;
  assign n1674 = ~n1468 & n1545;
  assign n1675 = n1471 & ~n1563;
  assign n1676 = ~n1471 & n1563;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = ~n1545 & n1677;
  assign n1679 = ~n1674 & ~n1678;
  assign n1680 = pi07 & ~n1679;
  assign n1681 = ~n1673 & n1680;
  assign n1682 = pi08 & ~n1672;
  assign n1683 = pi09 & ~n1665;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = ~n1681 & n1684;
  assign n1686 = ~n1659 & ~n1666;
  assign n1687 = ~n1685 & n1686;
  assign n1688 = ~n1658 & ~n1687;
  assign n1689 = n1651 & n1688;
  assign n1690 = ~n1648 & ~n1689;
  assign n1691 = ~n1525 & n1545;
  assign n1692 = ~n1528 & ~n1561;
  assign n1693 = n1528 & n1561;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = ~n1545 & n1694;
  assign n1696 = ~n1691 & ~n1695;
  assign n1697 = ~pi06 & n1696;
  assign n1698 = pi06 & ~n1696;
  assign n1699 = ~n1509 & n1545;
  assign n1700 = n1512 & ~n1559;
  assign n1701 = ~n1512 & n1559;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1545 & n1702;
  assign n1704 = ~n1699 & ~n1703;
  assign n1705 = ~pi05 & n1704;
  assign n1706 = ~n1500 & n1545;
  assign n1707 = n1503 & ~n1557;
  assign n1708 = ~n1503 & n1557;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1545 & n1709;
  assign n1711 = ~n1706 & ~n1710;
  assign n1712 = ~pi04 & n1711;
  assign n1713 = ~n1519 & ~n1541;
  assign n1714 = n1540 & ~n1713;
  assign n1715 = ~n1540 & n1713;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = ~n1545 & ~n1716;
  assign n1718 = n1518 & n1545;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = pi03 & n1719;
  assign n1721 = ~n1712 & n1720;
  assign n1722 = pi04 & ~n1711;
  assign n1723 = pi05 & ~n1704;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~n1721 & n1724;
  assign n1726 = ~n1705 & ~n1725;
  assign n1727 = ~n1698 & ~n1726;
  assign n1728 = ~n1658 & ~n1659;
  assign n1729 = ~n1673 & ~n1682;
  assign n1730 = ~pi07 & n1679;
  assign n1731 = ~n1680 & ~n1730;
  assign n1732 = ~n1666 & ~n1683;
  assign n1733 = n1729 & n1731;
  assign n1734 = n1732 & n1733;
  assign n1735 = n1728 & n1734;
  assign n1736 = n1651 & n1735;
  assign n1737 = ~n1697 & ~n1727;
  assign n1738 = n1736 & n1737;
  assign n1739 = ~n1690 & ~n1738;
  assign n1740 = ~n1697 & ~n1698;
  assign n1741 = ~n1712 & ~n1722;
  assign n1742 = ~pi03 & ~n1719;
  assign n1743 = ~n1720 & ~n1742;
  assign n1744 = ~n1705 & ~n1723;
  assign n1745 = n1740 & n1741;
  assign n1746 = n1743 & n1744;
  assign n1747 = n1745 & n1746;
  assign n1748 = n1736 & n1747;
  assign n1749 = ~n1739 & ~n1748;
  assign n1750 = pi02 & ~n1553;
  assign n1751 = ~pi02 & n1553;
  assign n1752 = pi00 & ~n1545;
  assign n1753 = ~pi01 & n1752;
  assign n1754 = ~n1751 & ~n1753;
  assign n1755 = ~n1750 & ~n1754;
  assign n1756 = n1748 & ~n1755;
  assign n1757 = ~n1749 & ~n1756;
  assign n1758 = ~n1750 & ~n1751;
  assign n1759 = n84 & n1758;
  assign n1760 = n1748 & n1759;
  assign n1761 = ~n1757 & ~n1760;
  assign n1762 = ~n1553 & n1761;
  assign n1763 = ~n84 & ~n1753;
  assign n1764 = ~n1758 & ~n1763;
  assign n1765 = n1758 & n1763;
  assign n1766 = ~n1764 & ~n1765;
  assign n1767 = ~n1761 & n1766;
  assign n1768 = ~n1762 & ~n1767;
  assign n1769 = n1576 & n1761;
  assign n1770 = ~n1751 & n1763;
  assign n1771 = ~n1750 & ~n1770;
  assign n1772 = ~n1720 & n1771;
  assign n1773 = ~n1742 & ~n1772;
  assign n1774 = ~n1712 & n1773;
  assign n1775 = ~n1722 & ~n1774;
  assign n1776 = ~n1723 & n1775;
  assign n1777 = ~n1705 & ~n1776;
  assign n1778 = ~n1697 & n1777;
  assign n1779 = ~n1698 & ~n1778;
  assign n1780 = ~n1730 & ~n1779;
  assign n1781 = ~n1680 & ~n1780;
  assign n1782 = ~n1673 & ~n1781;
  assign n1783 = ~n1682 & ~n1782;
  assign n1784 = ~n1683 & n1783;
  assign n1785 = ~n1666 & ~n1784;
  assign n1786 = ~n1659 & n1785;
  assign n1787 = ~n1658 & ~n1786;
  assign n1788 = n1650 & ~n1787;
  assign n1789 = ~n1650 & n1787;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1761 & n1790;
  assign n1792 = ~n1769 & ~n1791;
  assign n1793 = pi12 & ~n1792;
  assign n1794 = ~n1593 & n1761;
  assign n1795 = ~n1649 & n1787;
  assign n1796 = ~n1577 & ~n1795;
  assign n1797 = ~n1604 & n1796;
  assign n1798 = ~n1603 & ~n1797;
  assign n1799 = ~n1621 & n1798;
  assign n1800 = ~n1622 & ~n1799;
  assign n1801 = ~n1631 & n1800;
  assign n1802 = ~n1630 & ~n1801;
  assign n1803 = ~n1613 & ~n1802;
  assign n1804 = ~n1612 & ~n1803;
  assign n1805 = n1596 & ~n1804;
  assign n1806 = ~n1596 & n1804;
  assign n1807 = ~n1761 & ~n1805;
  assign n1808 = ~n1806 & n1807;
  assign n1809 = ~n1794 & ~n1808;
  assign n1810 = ~pi17 & n1809;
  assign n1811 = pi17 & ~n1809;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = ~n1611 & n1761;
  assign n1814 = n1614 & ~n1802;
  assign n1815 = ~n1614 & n1802;
  assign n1816 = ~n1761 & ~n1814;
  assign n1817 = ~n1815 & n1816;
  assign n1818 = ~n1813 & ~n1817;
  assign n1819 = ~pi16 & n1818;
  assign n1820 = pi16 & ~n1818;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = ~n1620 & n1761;
  assign n1823 = n1623 & ~n1798;
  assign n1824 = ~n1623 & n1798;
  assign n1825 = ~n1761 & ~n1823;
  assign n1826 = ~n1824 & n1825;
  assign n1827 = ~n1822 & ~n1826;
  assign n1828 = ~pi14 & n1827;
  assign n1829 = pi14 & ~n1827;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~n1602 & n1761;
  assign n1832 = ~n1605 & ~n1796;
  assign n1833 = n1605 & n1796;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = ~n1761 & n1834;
  assign n1836 = ~n1831 & ~n1835;
  assign n1837 = pi13 & ~n1836;
  assign n1838 = ~pi13 & n1836;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = ~pi12 & n1792;
  assign n1841 = ~n1629 & n1761;
  assign n1842 = ~n1632 & ~n1800;
  assign n1843 = n1632 & n1800;
  assign n1844 = ~n1761 & ~n1842;
  assign n1845 = ~n1843 & n1844;
  assign n1846 = ~n1841 & ~n1845;
  assign n1847 = pi15 & ~n1846;
  assign n1848 = ~pi15 & n1846;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = n1416 & ~n1840;
  assign n1851 = n1839 & n1850;
  assign n1852 = n1830 & n1851;
  assign n1853 = n1849 & n1852;
  assign n1854 = n1821 & n1853;
  assign n1855 = n1812 & n1854;
  assign n1856 = ~n1793 & n1855;
  assign n1857 = ~n1665 & n1761;
  assign n1858 = n1732 & ~n1783;
  assign n1859 = ~n1732 & n1783;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1761 & n1860;
  assign n1862 = ~n1857 & ~n1861;
  assign n1863 = ~pi10 & n1862;
  assign n1864 = pi10 & ~n1862;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1672 & n1761;
  assign n1867 = n1729 & ~n1781;
  assign n1868 = ~n1729 & n1781;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = ~n1761 & n1869;
  assign n1871 = ~n1866 & ~n1870;
  assign n1872 = pi09 & ~n1871;
  assign n1873 = ~pi09 & n1871;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1657 & n1761;
  assign n1876 = ~n1728 & ~n1785;
  assign n1877 = n1728 & n1785;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n1761 & n1878;
  assign n1880 = ~n1875 & ~n1879;
  assign n1881 = pi11 & ~n1880;
  assign n1882 = ~pi11 & n1880;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = ~n1679 & n1761;
  assign n1885 = n1731 & ~n1779;
  assign n1886 = ~n1731 & n1779;
  assign n1887 = ~n1885 & ~n1886;
  assign n1888 = ~n1761 & n1887;
  assign n1889 = ~n1884 & ~n1888;
  assign n1890 = pi08 & ~n1889;
  assign n1891 = ~pi08 & n1889;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = n1865 & n1874;
  assign n1894 = n1883 & n1892;
  assign n1895 = n1893 & n1894;
  assign n1896 = n1856 & n1895;
  assign n1897 = ~n1696 & n1761;
  assign n1898 = ~n1740 & ~n1777;
  assign n1899 = n1740 & n1777;
  assign n1900 = ~n1898 & ~n1899;
  assign n1901 = ~n1761 & n1900;
  assign n1902 = ~n1897 & ~n1901;
  assign n1903 = ~pi07 & n1902;
  assign n1904 = ~n1704 & n1761;
  assign n1905 = n1744 & ~n1775;
  assign n1906 = ~n1744 & n1775;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~n1761 & n1907;
  assign n1909 = ~n1904 & ~n1908;
  assign n1910 = pi06 & ~n1909;
  assign n1911 = pi07 & ~n1902;
  assign n1912 = ~pi06 & n1909;
  assign n1913 = ~n1711 & n1761;
  assign n1914 = ~n1741 & ~n1773;
  assign n1915 = n1741 & n1773;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = ~n1761 & n1916;
  assign n1918 = ~n1913 & ~n1917;
  assign n1919 = ~pi05 & n1918;
  assign n1920 = n1719 & n1761;
  assign n1921 = n1743 & ~n1771;
  assign n1922 = ~n1743 & n1771;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = ~n1761 & n1923;
  assign n1925 = ~n1920 & ~n1924;
  assign n1926 = ~pi04 & n1925;
  assign n1927 = pi05 & ~n1918;
  assign n1928 = n1926 & ~n1927;
  assign n1929 = ~n1912 & ~n1919;
  assign n1930 = ~n1928 & n1929;
  assign n1931 = ~n1910 & ~n1911;
  assign n1932 = ~n1930 & n1931;
  assign n1933 = ~n1903 & ~n1932;
  assign n1934 = n1896 & n1933;
  assign n1935 = ~n1872 & ~n1890;
  assign n1936 = ~n1863 & ~n1873;
  assign n1937 = ~n1935 & n1936;
  assign n1938 = ~n1864 & ~n1881;
  assign n1939 = ~n1937 & n1938;
  assign n1940 = ~n1882 & ~n1939;
  assign n1941 = n1856 & ~n1940;
  assign n1942 = ~n1829 & ~n1837;
  assign n1943 = ~n1828 & ~n1942;
  assign n1944 = ~n1848 & n1943;
  assign n1945 = ~n1847 & ~n1944;
  assign n1946 = ~n1820 & n1945;
  assign n1947 = ~n1819 & ~n1946;
  assign n1948 = ~n1810 & n1947;
  assign n1949 = n1416 & ~n1811;
  assign n1950 = ~n1948 & n1949;
  assign n1951 = ~n1855 & n1950;
  assign n1952 = ~n1941 & ~n1951;
  assign n1953 = ~n1934 & ~n1952;
  assign n1954 = ~n1919 & ~n1927;
  assign n1955 = pi04 & ~n1925;
  assign n1956 = ~n1926 & ~n1955;
  assign n1957 = ~n1903 & ~n1911;
  assign n1958 = ~n1910 & ~n1912;
  assign n1959 = n1954 & n1956;
  assign n1960 = n1957 & n1958;
  assign n1961 = n1959 & n1960;
  assign n1962 = n1896 & n1961;
  assign n1963 = ~pi03 & n1768;
  assign n1964 = pi03 & ~n1768;
  assign n1965 = pi00 & ~n1538;
  assign n1966 = n1543 & n1551;
  assign n1967 = ~pi01 & ~n1966;
  assign n1968 = n1965 & n1967;
  assign n1969 = pi01 & ~n1965;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~n1761 & n1970;
  assign n1972 = ~n1752 & n1761;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = pi02 & ~n1973;
  assign n1975 = ~n1964 & ~n1974;
  assign n1976 = ~n1963 & ~n1975;
  assign n1977 = n1962 & ~n1976;
  assign n1978 = ~n1953 & ~n1977;
  assign n1979 = ~pi02 & n1973;
  assign n1980 = ~n1974 & ~n1979;
  assign n1981 = ~n1963 & ~n1964;
  assign n1982 = n1980 & n1981;
  assign n1983 = n1962 & n1982;
  assign n1984 = ~n1978 & ~n1983;
  assign n1985 = pi00 & n1761;
  assign n1986 = ~pi01 & ~n1985;
  assign n1987 = n1983 & n1986;
  assign n1988 = ~n1984 & ~n1987;
  assign n1989 = ~n1768 & n1988;
  assign n1990 = ~n1979 & ~n1986;
  assign n1991 = ~n1974 & ~n1990;
  assign n1992 = n1981 & ~n1991;
  assign n1993 = ~n1981 & n1991;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = ~n1988 & n1994;
  assign n1996 = ~n1989 & ~n1995;
  assign n1997 = pi04 & ~n1996;
  assign n1998 = ~pi04 & n1996;
  assign n1999 = n1973 & n1988;
  assign n2000 = ~n1980 & ~n1986;
  assign n2001 = n1980 & n1986;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~n1988 & n2002;
  assign n2004 = ~n1999 & ~n2003;
  assign n2005 = pi03 & n2004;
  assign n2006 = pi00 & ~n1757;
  assign n2007 = ~pi01 & ~n2006;
  assign n2008 = pi01 & n2006;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n1988 & ~n2009;
  assign n2011 = pi00 & ~n1761;
  assign n2012 = n1988 & ~n2011;
  assign n2013 = ~n2010 & ~n2012;
  assign n2014 = ~pi02 & n2013;
  assign n2015 = pi02 & ~n2013;
  assign n2016 = pi00 & ~n1988;
  assign n2017 = ~pi01 & n2016;
  assign n2018 = ~n2015 & n2017;
  assign n2019 = ~pi03 & ~n2004;
  assign n2020 = ~n2014 & ~n2019;
  assign n2021 = ~n2018 & n2020;
  assign n2022 = ~n2005 & ~n2021;
  assign n2023 = ~n1998 & ~n2022;
  assign n2024 = n1792 & n1988;
  assign n2025 = ~n1793 & ~n1840;
  assign n2026 = ~n1964 & n1991;
  assign n2027 = ~n1963 & ~n2026;
  assign n2028 = ~n1955 & ~n2027;
  assign n2029 = ~n1926 & ~n2028;
  assign n2030 = ~n1927 & ~n2029;
  assign n2031 = ~n1919 & ~n2030;
  assign n2032 = ~n1912 & n2031;
  assign n2033 = ~n1910 & ~n2032;
  assign n2034 = ~n1903 & ~n2033;
  assign n2035 = ~n1911 & ~n2034;
  assign n2036 = ~n1891 & ~n2035;
  assign n2037 = ~n1890 & ~n2036;
  assign n2038 = ~n1872 & n2037;
  assign n2039 = ~n1873 & ~n2038;
  assign n2040 = ~n1864 & ~n2039;
  assign n2041 = ~n1863 & ~n2040;
  assign n2042 = ~n1882 & n2041;
  assign n2043 = ~n1881 & ~n2042;
  assign n2044 = ~n2025 & ~n2043;
  assign n2045 = n2025 & n2043;
  assign n2046 = ~n1988 & ~n2044;
  assign n2047 = ~n2045 & n2046;
  assign n2048 = ~n2024 & ~n2047;
  assign n2049 = pi13 & n2048;
  assign n2050 = ~pi13 & ~n2048;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = ~n1809 & n1988;
  assign n2053 = ~n1840 & ~n2043;
  assign n2054 = ~n1793 & ~n2053;
  assign n2055 = ~n1838 & ~n2054;
  assign n2056 = ~n1837 & ~n2055;
  assign n2057 = ~n1829 & n2056;
  assign n2058 = ~n1828 & ~n2057;
  assign n2059 = ~n1848 & n2058;
  assign n2060 = ~n1847 & ~n2059;
  assign n2061 = ~n1819 & ~n2060;
  assign n2062 = ~n1820 & ~n2061;
  assign n2063 = n1812 & ~n2062;
  assign n2064 = ~n1812 & n2062;
  assign n2065 = ~n1988 & ~n2063;
  assign n2066 = ~n2064 & n2065;
  assign n2067 = ~n2052 & ~n2066;
  assign n2068 = pi18 & ~n2067;
  assign n2069 = ~pi18 & n2067;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n1846 & n1988;
  assign n2072 = ~n1849 & ~n2058;
  assign n2073 = n1849 & n2058;
  assign n2074 = ~n1988 & ~n2072;
  assign n2075 = ~n2073 & n2074;
  assign n2076 = ~n2071 & ~n2075;
  assign n2077 = pi16 & ~n2076;
  assign n2078 = ~pi16 & n2076;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = ~n1818 & n1988;
  assign n2081 = n1821 & ~n2060;
  assign n2082 = ~n1821 & n2060;
  assign n2083 = ~n1988 & ~n2081;
  assign n2084 = ~n2082 & n2083;
  assign n2085 = ~n2080 & ~n2084;
  assign n2086 = pi17 & ~n2085;
  assign n2087 = ~pi17 & n2085;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = ~n1827 & n1988;
  assign n2090 = n1830 & ~n2056;
  assign n2091 = ~n1830 & n2056;
  assign n2092 = ~n1988 & ~n2090;
  assign n2093 = ~n2091 & n2092;
  assign n2094 = ~n2089 & ~n2093;
  assign n2095 = pi15 & ~n2094;
  assign n2096 = ~pi15 & n2094;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = ~n1836 & n1988;
  assign n2099 = n1839 & ~n2054;
  assign n2100 = ~n1839 & n2054;
  assign n2101 = ~n1988 & ~n2099;
  assign n2102 = ~n2100 & n2101;
  assign n2103 = ~n2098 & ~n2102;
  assign n2104 = pi14 & ~n2103;
  assign n2105 = ~pi14 & n2103;
  assign n2106 = ~n2104 & ~n2105;
  assign n2107 = n76 & n2106;
  assign n2108 = n2097 & n2107;
  assign n2109 = n2079 & n2108;
  assign n2110 = n2088 & n2109;
  assign n2111 = n2070 & n2110;
  assign n2112 = n2051 & n2111;
  assign n2113 = n1880 & n1988;
  assign n2114 = n1883 & ~n2041;
  assign n2115 = ~n1883 & n2041;
  assign n2116 = ~n1988 & ~n2114;
  assign n2117 = ~n2115 & n2116;
  assign n2118 = ~n2113 & ~n2117;
  assign n2119 = pi12 & n2118;
  assign n2120 = ~pi12 & ~n2118;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = ~n1889 & n1988;
  assign n2123 = n1892 & ~n2035;
  assign n2124 = ~n1892 & n2035;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = ~n1988 & n2125;
  assign n2127 = ~n2122 & ~n2126;
  assign n2128 = pi09 & ~n2127;
  assign n2129 = ~pi09 & n2127;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n1871 & n1988;
  assign n2132 = n1874 & ~n2037;
  assign n2133 = ~n1874 & n2037;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = ~n1988 & n2134;
  assign n2136 = ~n2131 & ~n2135;
  assign n2137 = pi10 & ~n2136;
  assign n2138 = ~pi10 & n2136;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = n1862 & n1988;
  assign n2141 = n1865 & ~n2039;
  assign n2142 = ~n1865 & n2039;
  assign n2143 = ~n1988 & ~n2141;
  assign n2144 = ~n2142 & n2143;
  assign n2145 = ~n2140 & ~n2144;
  assign n2146 = pi11 & n2145;
  assign n2147 = ~pi11 & ~n2145;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = n2130 & n2139;
  assign n2150 = n2148 & n2149;
  assign n2151 = n2121 & n2150;
  assign n2152 = n2112 & n2151;
  assign n2153 = ~n1909 & n1988;
  assign n2154 = ~n1958 & ~n2031;
  assign n2155 = n1958 & n2031;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~n1988 & n2156;
  assign n2158 = ~n2153 & ~n2157;
  assign n2159 = pi07 & ~n2158;
  assign n2160 = ~pi07 & n2158;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~n1918 & n1988;
  assign n2163 = ~n1954 & ~n2029;
  assign n2164 = n1954 & n2029;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = ~n1988 & n2165;
  assign n2167 = ~n2162 & ~n2166;
  assign n2168 = pi06 & ~n2167;
  assign n2169 = ~pi06 & n2167;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = ~n1925 & n1988;
  assign n2172 = ~n1956 & ~n2027;
  assign n2173 = n1956 & n2027;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175 = ~n1988 & n2174;
  assign n2176 = ~n2171 & ~n2175;
  assign n2177 = pi05 & ~n2176;
  assign n2178 = ~pi05 & n2176;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n1902 & n1988;
  assign n2181 = n1957 & ~n2033;
  assign n2182 = ~n1957 & n2033;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = ~n1988 & n2183;
  assign n2185 = ~n2180 & ~n2184;
  assign n2186 = pi08 & ~n2185;
  assign n2187 = ~pi08 & n2185;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = n2161 & n2170;
  assign n2190 = n2179 & n2188;
  assign n2191 = n2189 & n2190;
  assign n2192 = n2152 & n2191;
  assign n2193 = ~n1997 & ~n2023;
  assign n2194 = n2192 & n2193;
  assign n2195 = ~n2050 & n2111;
  assign n2196 = ~n2095 & ~n2104;
  assign n2197 = ~n2096 & ~n2196;
  assign n2198 = ~n2078 & n2197;
  assign n2199 = ~n2077 & ~n2198;
  assign n2200 = ~n2086 & n2199;
  assign n2201 = ~n2087 & ~n2200;
  assign n2202 = ~n2069 & n2201;
  assign n2203 = n76 & ~n2068;
  assign n2204 = ~n2202 & n2203;
  assign n2205 = ~n2195 & n2204;
  assign n2206 = ~n2128 & ~n2137;
  assign n2207 = ~n2138 & ~n2147;
  assign n2208 = ~n2206 & n2207;
  assign n2209 = ~n2119 & ~n2146;
  assign n2210 = ~n2208 & n2209;
  assign n2211 = ~n2120 & ~n2210;
  assign n2212 = n2112 & ~n2211;
  assign n2213 = ~n2205 & ~n2212;
  assign n2214 = ~n2169 & ~n2178;
  assign n2215 = ~n2159 & ~n2168;
  assign n2216 = ~n2214 & n2215;
  assign n2217 = ~n2160 & ~n2187;
  assign n2218 = ~n2216 & n2217;
  assign n2219 = ~n2186 & ~n2218;
  assign n2220 = n2152 & ~n2219;
  assign n2221 = ~n2213 & ~n2220;
  assign n2222 = ~n2194 & ~n2221;
  assign n2223 = ~n2014 & ~n2015;
  assign n2224 = ~n1997 & ~n1998;
  assign n2225 = ~n2005 & ~n2019;
  assign n2226 = n84 & n2223;
  assign n2227 = n2224 & n2225;
  assign n2228 = n2226 & n2227;
  assign n2229 = n2192 & n2228;
  assign n2230 = n2222 & ~n2229;
  assign n2231 = pi00 & ~n2230;
  assign n2232 = ~pi01 & n2231;
  assign n2233 = ~n2176 & n2230;
  assign n2234 = ~n84 & ~n2017;
  assign n2235 = ~n2014 & n2234;
  assign n2236 = ~n2015 & ~n2235;
  assign n2237 = ~n2019 & ~n2236;
  assign n2238 = ~n2005 & ~n2237;
  assign n2239 = ~n1998 & ~n2238;
  assign n2240 = ~n1997 & ~n2239;
  assign n2241 = n2179 & ~n2240;
  assign n2242 = ~n2179 & n2240;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = ~n2230 & n2243;
  assign n2245 = ~n2233 & ~n2244;
  assign n2246 = pi06 & ~n2245;
  assign n2247 = ~n2118 & n2230;
  assign n2248 = ~n2178 & ~n2240;
  assign n2249 = ~n2177 & ~n2248;
  assign n2250 = ~n2169 & ~n2249;
  assign n2251 = ~n2168 & ~n2250;
  assign n2252 = ~n2160 & ~n2251;
  assign n2253 = ~n2159 & ~n2252;
  assign n2254 = ~n2186 & n2253;
  assign n2255 = ~n2187 & ~n2254;
  assign n2256 = ~n2128 & ~n2255;
  assign n2257 = ~n2129 & ~n2256;
  assign n2258 = ~n2138 & n2257;
  assign n2259 = ~n2137 & ~n2258;
  assign n2260 = ~n2146 & n2259;
  assign n2261 = ~n2147 & ~n2260;
  assign n2262 = n2121 & ~n2261;
  assign n2263 = ~n2121 & n2261;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = ~n2230 & n2264;
  assign n2266 = ~n2247 & ~n2265;
  assign n2267 = pi13 & n2266;
  assign n2268 = ~pi13 & ~n2266;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = n2145 & n2230;
  assign n2271 = n2148 & ~n2259;
  assign n2272 = ~n2148 & n2259;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = ~n2230 & n2273;
  assign n2275 = ~n2270 & ~n2274;
  assign n2276 = pi12 & ~n2275;
  assign n2277 = ~pi12 & n2275;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~n2130 & ~n2255;
  assign n2280 = n2130 & n2255;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = ~n2230 & ~n2281;
  assign n2283 = n2127 & n2230;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = pi10 & n2284;
  assign n2286 = ~pi10 & ~n2284;
  assign n2287 = ~n2285 & ~n2286;
  assign n2288 = ~n2048 & n2230;
  assign n2289 = ~n2119 & ~n2261;
  assign n2290 = ~n2120 & ~n2289;
  assign n2291 = n2051 & ~n2290;
  assign n2292 = ~n2051 & n2290;
  assign n2293 = ~n2230 & ~n2291;
  assign n2294 = ~n2292 & n2293;
  assign n2295 = ~n2288 & ~n2294;
  assign n2296 = pi14 & n2295;
  assign n2297 = ~n2103 & n2230;
  assign n2298 = ~n2049 & ~n2290;
  assign n2299 = ~n2050 & ~n2298;
  assign n2300 = ~n2106 & ~n2299;
  assign n2301 = n2106 & n2299;
  assign n2302 = ~n2230 & ~n2300;
  assign n2303 = ~n2301 & n2302;
  assign n2304 = ~n2297 & ~n2303;
  assign n2305 = pi15 & ~n2304;
  assign n2306 = ~pi15 & n2304;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n2076 & n2230;
  assign n2309 = ~n2105 & n2299;
  assign n2310 = ~n2104 & ~n2309;
  assign n2311 = ~n2095 & n2310;
  assign n2312 = ~n2096 & ~n2311;
  assign n2313 = ~n2079 & ~n2312;
  assign n2314 = n2079 & n2312;
  assign n2315 = ~n2230 & ~n2313;
  assign n2316 = ~n2314 & n2315;
  assign n2317 = ~n2308 & ~n2316;
  assign n2318 = pi17 & ~n2317;
  assign n2319 = ~pi17 & n2317;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~pi14 & ~n2295;
  assign n2322 = ~pi20 & n75;
  assign n2323 = ~n2094 & n2230;
  assign n2324 = n2097 & ~n2310;
  assign n2325 = ~n2097 & n2310;
  assign n2326 = ~n2230 & ~n2324;
  assign n2327 = ~n2325 & n2326;
  assign n2328 = ~n2323 & ~n2327;
  assign n2329 = pi16 & ~n2328;
  assign n2330 = ~pi16 & n2328;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = ~n2067 & n2230;
  assign n2333 = ~n2078 & n2312;
  assign n2334 = ~n2077 & ~n2333;
  assign n2335 = ~n2087 & ~n2334;
  assign n2336 = ~n2086 & ~n2335;
  assign n2337 = n2070 & ~n2336;
  assign n2338 = ~n2070 & n2336;
  assign n2339 = ~n2230 & ~n2337;
  assign n2340 = ~n2338 & n2339;
  assign n2341 = ~n2332 & ~n2340;
  assign n2342 = pi19 & ~n2341;
  assign n2343 = ~pi19 & n2341;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = ~n2085 & n2230;
  assign n2346 = n2088 & ~n2334;
  assign n2347 = ~n2088 & n2334;
  assign n2348 = ~n2230 & ~n2346;
  assign n2349 = ~n2347 & n2348;
  assign n2350 = ~n2345 & ~n2349;
  assign n2351 = pi18 & ~n2350;
  assign n2352 = ~pi18 & n2350;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~n2321 & n2322;
  assign n2355 = n2307 & n2354;
  assign n2356 = n2331 & n2355;
  assign n2357 = n2320 & n2356;
  assign n2358 = n2353 & n2357;
  assign n2359 = n2344 & n2358;
  assign n2360 = ~n2296 & n2359;
  assign n2361 = ~n2136 & n2230;
  assign n2362 = ~n2139 & ~n2257;
  assign n2363 = n2139 & n2257;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = ~n2230 & n2364;
  assign n2366 = ~n2361 & ~n2365;
  assign n2367 = pi11 & ~n2366;
  assign n2368 = ~pi11 & n2366;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = n2269 & n2278;
  assign n2371 = n2287 & n2369;
  assign n2372 = n2370 & n2371;
  assign n2373 = n2360 & n2372;
  assign n2374 = ~n2167 & n2230;
  assign n2375 = n2170 & ~n2249;
  assign n2376 = ~n2170 & n2249;
  assign n2377 = ~n2375 & ~n2376;
  assign n2378 = ~n2230 & n2377;
  assign n2379 = ~n2374 & ~n2378;
  assign n2380 = pi07 & ~n2379;
  assign n2381 = ~pi07 & n2379;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = ~n2185 & n2230;
  assign n2384 = n2188 & ~n2253;
  assign n2385 = ~n2188 & n2253;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~n2230 & n2386;
  assign n2388 = ~n2383 & ~n2387;
  assign n2389 = pi09 & ~n2388;
  assign n2390 = ~pi09 & n2388;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = ~pi06 & n2245;
  assign n2393 = n2158 & n2230;
  assign n2394 = ~n2161 & ~n2251;
  assign n2395 = n2161 & n2251;
  assign n2396 = ~n2394 & ~n2395;
  assign n2397 = ~n2230 & n2396;
  assign n2398 = ~n2393 & ~n2397;
  assign n2399 = pi08 & n2398;
  assign n2400 = ~pi08 & ~n2398;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = n2382 & ~n2392;
  assign n2403 = n2391 & n2401;
  assign n2404 = n2402 & n2403;
  assign n2405 = ~n2246 & n2404;
  assign n2406 = n2373 & n2405;
  assign n2407 = ~n1996 & n2230;
  assign n2408 = n2224 & ~n2238;
  assign n2409 = ~n2224 & n2238;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n2230 & n2410;
  assign n2412 = ~n2407 & ~n2411;
  assign n2413 = pi05 & ~n2412;
  assign n2414 = ~pi05 & n2412;
  assign n2415 = ~n2413 & ~n2414;
  assign n2416 = n2004 & n2230;
  assign n2417 = n2225 & ~n2236;
  assign n2418 = ~n2225 & n2236;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = ~n2230 & n2419;
  assign n2421 = ~n2416 & ~n2420;
  assign n2422 = pi04 & ~n2421;
  assign n2423 = ~pi04 & n2421;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2013 & n2230;
  assign n2426 = ~n2223 & ~n2234;
  assign n2427 = n2223 & n2234;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n2230 & n2428;
  assign n2430 = ~n2425 & ~n2429;
  assign n2431 = ~pi03 & n2430;
  assign n2432 = pi03 & ~n2430;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = pi00 & ~n1984;
  assign n2435 = n1983 & n2011;
  assign n2436 = ~pi01 & ~n2435;
  assign n2437 = n2434 & n2436;
  assign n2438 = pi01 & ~n2434;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = ~n2230 & n2439;
  assign n2441 = ~n2016 & n2230;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = pi02 & ~n2442;
  assign n2444 = ~pi02 & n2442;
  assign n2445 = ~n2443 & ~n2444;
  assign n2446 = n2415 & n2424;
  assign n2447 = n2433 & n2445;
  assign n2448 = n2446 & n2447;
  assign n2449 = n2406 & n2448;
  assign n2450 = ~n2232 & n2449;
  assign n2451 = ~n2432 & ~n2443;
  assign n2452 = ~n2423 & ~n2431;
  assign n2453 = ~n2451 & n2452;
  assign n2454 = ~n2413 & ~n2422;
  assign n2455 = ~n2453 & n2454;
  assign n2456 = ~n2414 & ~n2455;
  assign n2457 = n2406 & ~n2456;
  assign n2458 = n2305 & ~n2330;
  assign n2459 = ~n2329 & ~n2458;
  assign n2460 = ~n2319 & ~n2459;
  assign n2461 = ~n2318 & ~n2460;
  assign n2462 = ~n2352 & ~n2461;
  assign n2463 = ~n2351 & ~n2462;
  assign n2464 = ~n2342 & n2463;
  assign n2465 = ~n2343 & ~n2464;
  assign n2466 = n2322 & ~n2359;
  assign n2467 = ~n2465 & n2466;
  assign n2468 = n2285 & ~n2368;
  assign n2469 = ~n2276 & ~n2367;
  assign n2470 = ~n2468 & n2469;
  assign n2471 = ~n2268 & ~n2277;
  assign n2472 = ~n2470 & n2471;
  assign n2473 = ~n2267 & ~n2472;
  assign n2474 = n2360 & n2473;
  assign n2475 = ~n2373 & ~n2467;
  assign n2476 = ~n2474 & n2475;
  assign n2477 = ~n2380 & ~n2399;
  assign n2478 = ~n2390 & ~n2400;
  assign n2479 = ~n2477 & n2478;
  assign n2480 = ~n2389 & ~n2479;
  assign n2481 = ~n2404 & n2480;
  assign n2482 = n2373 & ~n2481;
  assign n2483 = ~n2476 & ~n2482;
  assign n2484 = ~n2457 & ~n2483;
  assign n2485 = ~n2450 & ~n2484;
  assign n2486 = pi00 & n2485;
  assign n2487 = n84 & n2449;
  assign n2488 = ~n2485 & ~n2487;
  assign n2489 = n2295 & n2488;
  assign n2490 = ~n84 & ~n2232;
  assign n2491 = ~n2443 & ~n2490;
  assign n2492 = ~n2444 & ~n2491;
  assign n2493 = ~n2431 & n2492;
  assign n2494 = ~n2432 & ~n2493;
  assign n2495 = ~n2423 & ~n2494;
  assign n2496 = ~n2422 & ~n2495;
  assign n2497 = ~n2414 & ~n2496;
  assign n2498 = ~n2413 & ~n2497;
  assign n2499 = ~n2392 & ~n2498;
  assign n2500 = ~n2246 & ~n2499;
  assign n2501 = ~n2381 & ~n2500;
  assign n2502 = ~n2380 & ~n2501;
  assign n2503 = ~n2399 & n2502;
  assign n2504 = ~n2400 & ~n2503;
  assign n2505 = ~n2389 & ~n2504;
  assign n2506 = ~n2390 & ~n2505;
  assign n2507 = ~n2285 & ~n2506;
  assign n2508 = ~n2286 & ~n2507;
  assign n2509 = ~n2368 & n2508;
  assign n2510 = ~n2367 & ~n2509;
  assign n2511 = ~n2276 & n2510;
  assign n2512 = ~n2277 & ~n2511;
  assign n2513 = ~n2267 & ~n2512;
  assign n2514 = ~n2268 & ~n2513;
  assign n2515 = ~n2296 & ~n2321;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = n2514 & n2515;
  assign n2518 = ~n2488 & ~n2516;
  assign n2519 = ~n2517 & n2518;
  assign n2520 = ~n2489 & ~n2519;
  assign n2521 = ~pi15 & n2520;
  assign n2522 = ~n2341 & n2488;
  assign n2523 = ~n2296 & ~n2514;
  assign n2524 = ~n2321 & ~n2523;
  assign n2525 = ~n2305 & ~n2524;
  assign n2526 = ~n2306 & ~n2525;
  assign n2527 = ~n2330 & n2526;
  assign n2528 = ~n2329 & ~n2527;
  assign n2529 = ~n2319 & ~n2528;
  assign n2530 = ~n2318 & ~n2529;
  assign n2531 = ~n2352 & ~n2530;
  assign n2532 = ~n2351 & ~n2531;
  assign n2533 = n2344 & ~n2532;
  assign n2534 = ~n2344 & n2532;
  assign n2535 = ~n2488 & ~n2533;
  assign n2536 = ~n2534 & n2535;
  assign n2537 = ~n2522 & ~n2536;
  assign n2538 = pi20 & ~n2537;
  assign n2539 = ~pi20 & n2537;
  assign n2540 = ~n2538 & ~n2539;
  assign n2541 = ~n2317 & n2488;
  assign n2542 = n2320 & ~n2528;
  assign n2543 = ~n2320 & n2528;
  assign n2544 = ~n2488 & ~n2542;
  assign n2545 = ~n2543 & n2544;
  assign n2546 = ~n2541 & ~n2545;
  assign n2547 = pi18 & ~n2546;
  assign n2548 = ~pi18 & n2546;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = ~n2350 & n2488;
  assign n2551 = n2353 & ~n2530;
  assign n2552 = ~n2353 & n2530;
  assign n2553 = ~n2488 & ~n2551;
  assign n2554 = ~n2552 & n2553;
  assign n2555 = ~n2550 & ~n2554;
  assign n2556 = pi19 & ~n2555;
  assign n2557 = ~pi19 & n2555;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = ~n2328 & n2488;
  assign n2560 = ~n2331 & ~n2526;
  assign n2561 = n2331 & n2526;
  assign n2562 = ~n2488 & ~n2560;
  assign n2563 = ~n2561 & n2562;
  assign n2564 = ~n2559 & ~n2563;
  assign n2565 = pi17 & ~n2564;
  assign n2566 = ~pi17 & n2564;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = n2304 & n2488;
  assign n2569 = n2307 & ~n2524;
  assign n2570 = ~n2307 & n2524;
  assign n2571 = ~n2488 & ~n2569;
  assign n2572 = ~n2570 & n2571;
  assign n2573 = ~n2568 & ~n2572;
  assign n2574 = pi16 & n2573;
  assign n2575 = ~pi16 & ~n2573;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = n75 & n2576;
  assign n2578 = n2567 & n2577;
  assign n2579 = n2549 & n2578;
  assign n2580 = n2558 & n2579;
  assign n2581 = n2540 & n2580;
  assign n2582 = ~n2521 & n2581;
  assign n2583 = ~n2565 & ~n2574;
  assign n2584 = ~n2566 & ~n2583;
  assign n2585 = ~n2548 & n2584;
  assign n2586 = ~n2547 & ~n2585;
  assign n2587 = ~n2556 & n2586;
  assign n2588 = ~n2557 & ~n2587;
  assign n2589 = ~n2539 & n2588;
  assign n2590 = n75 & ~n2538;
  assign n2591 = ~n2589 & n2590;
  assign n2592 = ~n2582 & n2591;
  assign n2593 = pi15 & ~n2520;
  assign n2594 = ~n2521 & ~n2593;
  assign n2595 = n2581 & n2594;
  assign n2596 = ~n2266 & n2488;
  assign n2597 = n2269 & ~n2512;
  assign n2598 = ~n2269 & n2512;
  assign n2599 = ~n2488 & ~n2597;
  assign n2600 = ~n2598 & n2599;
  assign n2601 = ~n2596 & ~n2600;
  assign n2602 = ~pi14 & ~n2601;
  assign n2603 = pi14 & n2601;
  assign n2604 = ~n2275 & n2488;
  assign n2605 = n2278 & ~n2510;
  assign n2606 = ~n2278 & n2510;
  assign n2607 = ~n2488 & ~n2605;
  assign n2608 = ~n2606 & n2607;
  assign n2609 = ~n2604 & ~n2608;
  assign n2610 = pi13 & ~n2609;
  assign n2611 = ~pi13 & n2609;
  assign n2612 = n2366 & n2488;
  assign n2613 = n2369 & ~n2508;
  assign n2614 = ~n2369 & n2508;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = ~n2488 & n2615;
  assign n2617 = ~n2612 & ~n2616;
  assign n2618 = ~pi12 & ~n2617;
  assign n2619 = ~n2284 & n2488;
  assign n2620 = n2287 & ~n2506;
  assign n2621 = ~n2287 & n2506;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = ~n2488 & n2622;
  assign n2624 = ~n2619 & ~n2623;
  assign n2625 = pi11 & n2624;
  assign n2626 = pi12 & n2617;
  assign n2627 = ~n2625 & ~n2626;
  assign n2628 = ~n2611 & ~n2618;
  assign n2629 = ~n2627 & n2628;
  assign n2630 = ~n2603 & ~n2610;
  assign n2631 = ~n2629 & n2630;
  assign n2632 = ~n2602 & ~n2631;
  assign n2633 = n2595 & ~n2632;
  assign n2634 = ~n2592 & ~n2633;
  assign n2635 = n2388 & n2488;
  assign n2636 = n2391 & ~n2504;
  assign n2637 = ~n2391 & n2504;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = ~n2488 & n2638;
  assign n2640 = ~n2635 & ~n2639;
  assign n2641 = pi10 & n2640;
  assign n2642 = ~pi10 & ~n2640;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = ~n2379 & n2488;
  assign n2645 = n2382 & ~n2500;
  assign n2646 = ~n2382 & n2500;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = ~n2488 & n2647;
  assign n2649 = ~n2644 & ~n2648;
  assign n2650 = pi08 & ~n2649;
  assign n2651 = ~pi08 & n2649;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = ~n2246 & ~n2392;
  assign n2654 = ~n2498 & ~n2653;
  assign n2655 = n2498 & n2653;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = ~n2488 & ~n2656;
  assign n2658 = ~n2245 & n2488;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = ~pi07 & n2659;
  assign n2661 = n2398 & n2488;
  assign n2662 = n2401 & ~n2502;
  assign n2663 = ~n2401 & n2502;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = ~n2488 & n2664;
  assign n2666 = ~n2661 & ~n2665;
  assign n2667 = pi09 & ~n2666;
  assign n2668 = ~pi09 & n2666;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = n2643 & ~n2660;
  assign n2671 = n2652 & n2669;
  assign n2672 = n2670 & n2671;
  assign n2673 = n2650 & ~n2668;
  assign n2674 = ~n2641 & ~n2667;
  assign n2675 = ~n2673 & n2674;
  assign n2676 = ~n2642 & ~n2675;
  assign n2677 = ~n2672 & ~n2676;
  assign n2678 = ~n2602 & ~n2603;
  assign n2679 = ~pi11 & ~n2624;
  assign n2680 = ~n2625 & ~n2679;
  assign n2681 = ~n2618 & ~n2626;
  assign n2682 = ~n2610 & ~n2611;
  assign n2683 = n2680 & n2681;
  assign n2684 = n2682 & n2683;
  assign n2685 = n2678 & n2684;
  assign n2686 = n2595 & n2685;
  assign n2687 = ~n2677 & n2686;
  assign n2688 = ~n2634 & ~n2687;
  assign n2689 = pi07 & ~n2659;
  assign n2690 = n2672 & ~n2689;
  assign n2691 = n2686 & n2690;
  assign n2692 = n2412 & n2488;
  assign n2693 = ~n2415 & ~n2496;
  assign n2694 = n2415 & n2496;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = ~n2488 & n2695;
  assign n2697 = ~n2692 & ~n2696;
  assign n2698 = pi06 & n2697;
  assign n2699 = ~pi06 & ~n2697;
  assign n2700 = ~n2421 & n2488;
  assign n2701 = n2424 & ~n2494;
  assign n2702 = ~n2424 & n2494;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = ~n2488 & n2703;
  assign n2705 = ~n2700 & ~n2704;
  assign n2706 = ~pi05 & n2705;
  assign n2707 = ~n2430 & n2488;
  assign n2708 = ~n2433 & ~n2492;
  assign n2709 = n2433 & n2492;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = ~n2488 & n2710;
  assign n2712 = ~n2707 & ~n2711;
  assign n2713 = pi04 & ~n2712;
  assign n2714 = pi05 & ~n2705;
  assign n2715 = ~pi04 & n2712;
  assign n2716 = ~n2445 & ~n2490;
  assign n2717 = n2445 & n2490;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = ~n2488 & ~n2718;
  assign n2720 = n2442 & n2488;
  assign n2721 = ~n2719 & ~n2720;
  assign n2722 = pi03 & n2721;
  assign n2723 = ~n2715 & n2722;
  assign n2724 = ~n2713 & ~n2714;
  assign n2725 = ~n2723 & n2724;
  assign n2726 = ~n2699 & ~n2706;
  assign n2727 = ~n2725 & n2726;
  assign n2728 = ~n2698 & ~n2727;
  assign n2729 = n2691 & n2728;
  assign n2730 = ~n2688 & ~n2729;
  assign n2731 = n314 & n2222;
  assign n2732 = pi01 & ~n2222;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = ~n2488 & n2733;
  assign n2735 = ~n2231 & n2488;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = pi02 & ~n2736;
  assign n2738 = ~pi02 & n2736;
  assign n2739 = ~pi01 & n2486;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = ~n2737 & ~n2740;
  assign n2742 = ~n2713 & ~n2715;
  assign n2743 = ~n2698 & ~n2699;
  assign n2744 = ~n2706 & ~n2714;
  assign n2745 = ~pi03 & ~n2721;
  assign n2746 = ~n2722 & ~n2745;
  assign n2747 = n2742 & n2743;
  assign n2748 = n2744 & n2746;
  assign n2749 = n2747 & n2748;
  assign n2750 = n2691 & n2749;
  assign n2751 = ~n2741 & n2750;
  assign n2752 = ~n2730 & ~n2751;
  assign n2753 = ~n2737 & ~n2738;
  assign n2754 = n84 & n2753;
  assign n2755 = n2750 & n2754;
  assign n2756 = ~n2752 & ~n2755;
  assign n2757 = ~n2486 & n2756;
  assign n2758 = pi00 & ~n2485;
  assign n2759 = ~pi01 & ~n2758;
  assign n2760 = pi01 & n2758;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = ~n2756 & ~n2761;
  assign n2763 = ~n2757 & ~n2762;
  assign n2764 = ~n2660 & ~n2689;
  assign n2765 = ~n2738 & ~n2759;
  assign n2766 = ~n2737 & ~n2765;
  assign n2767 = ~n2722 & n2766;
  assign n2768 = ~n2745 & ~n2767;
  assign n2769 = ~n2715 & n2768;
  assign n2770 = ~n2713 & ~n2769;
  assign n2771 = ~n2706 & ~n2770;
  assign n2772 = ~n2714 & ~n2771;
  assign n2773 = ~n2699 & ~n2772;
  assign n2774 = ~n2698 & ~n2773;
  assign n2775 = ~n2764 & ~n2774;
  assign n2776 = n2764 & n2774;
  assign n2777 = ~n2775 & ~n2776;
  assign n2778 = ~n2756 & ~n2777;
  assign n2779 = ~n2659 & n2756;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = pi08 & ~n2780;
  assign n2782 = n2520 & n2756;
  assign n2783 = ~n2660 & ~n2774;
  assign n2784 = ~n2689 & ~n2783;
  assign n2785 = ~n2651 & ~n2784;
  assign n2786 = ~n2650 & ~n2785;
  assign n2787 = ~n2668 & ~n2786;
  assign n2788 = ~n2667 & ~n2787;
  assign n2789 = ~n2641 & n2788;
  assign n2790 = ~n2642 & ~n2789;
  assign n2791 = ~n2625 & ~n2790;
  assign n2792 = ~n2679 & ~n2791;
  assign n2793 = ~n2626 & ~n2792;
  assign n2794 = ~n2618 & ~n2793;
  assign n2795 = ~n2610 & ~n2794;
  assign n2796 = ~n2611 & ~n2795;
  assign n2797 = ~n2603 & ~n2796;
  assign n2798 = ~n2602 & ~n2797;
  assign n2799 = n2594 & ~n2798;
  assign n2800 = ~n2594 & n2798;
  assign n2801 = ~n2756 & ~n2799;
  assign n2802 = ~n2800 & n2801;
  assign n2803 = ~n2782 & ~n2802;
  assign n2804 = pi16 & n2803;
  assign n2805 = ~n2537 & n2756;
  assign n2806 = ~n2521 & n2798;
  assign n2807 = ~n2593 & ~n2806;
  assign n2808 = ~n2575 & ~n2807;
  assign n2809 = ~n2574 & ~n2808;
  assign n2810 = ~n2565 & n2809;
  assign n2811 = ~n2566 & ~n2810;
  assign n2812 = ~n2548 & n2811;
  assign n2813 = ~n2547 & ~n2812;
  assign n2814 = ~n2557 & ~n2813;
  assign n2815 = ~n2556 & ~n2814;
  assign n2816 = n2540 & ~n2815;
  assign n2817 = ~n2540 & n2815;
  assign n2818 = ~n2756 & ~n2816;
  assign n2819 = ~n2817 & n2818;
  assign n2820 = ~n2805 & ~n2819;
  assign n2821 = pi21 & ~n2820;
  assign n2822 = ~pi21 & n2820;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = ~n2555 & n2756;
  assign n2825 = n2558 & ~n2813;
  assign n2826 = ~n2558 & n2813;
  assign n2827 = ~n2756 & ~n2825;
  assign n2828 = ~n2826 & n2827;
  assign n2829 = ~n2824 & ~n2828;
  assign n2830 = pi20 & ~n2829;
  assign n2831 = ~pi20 & n2829;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n2564 & n2756;
  assign n2834 = ~n2567 & ~n2809;
  assign n2835 = n2567 & n2809;
  assign n2836 = ~n2756 & ~n2834;
  assign n2837 = ~n2835 & n2836;
  assign n2838 = ~n2833 & ~n2837;
  assign n2839 = pi18 & n2838;
  assign n2840 = ~pi18 & ~n2838;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2576 & ~n2807;
  assign n2843 = n2576 & n2807;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = ~n2756 & ~n2844;
  assign n2846 = n2573 & n2756;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = pi17 & ~n2847;
  assign n2849 = ~pi17 & n2847;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~pi16 & ~n2803;
  assign n2852 = ~n2546 & n2756;
  assign n2853 = ~n2549 & ~n2811;
  assign n2854 = n2549 & n2811;
  assign n2855 = ~n2756 & ~n2853;
  assign n2856 = ~n2854 & n2855;
  assign n2857 = ~n2852 & ~n2856;
  assign n2858 = pi19 & ~n2857;
  assign n2859 = ~pi19 & n2857;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = n74 & ~n2851;
  assign n2862 = n2850 & n2861;
  assign n2863 = n2841 & n2862;
  assign n2864 = n2860 & n2863;
  assign n2865 = n2832 & n2864;
  assign n2866 = n2823 & n2865;
  assign n2867 = ~n2804 & n2866;
  assign n2868 = ~n2678 & ~n2796;
  assign n2869 = n2678 & n2796;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = ~n2756 & ~n2870;
  assign n2872 = ~n2601 & n2756;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = pi15 & n2873;
  assign n2875 = ~pi15 & ~n2873;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = ~n2617 & n2756;
  assign n2878 = n2681 & ~n2792;
  assign n2879 = ~n2681 & n2792;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = ~n2756 & n2880;
  assign n2882 = ~n2877 & ~n2881;
  assign n2883 = pi13 & n2882;
  assign n2884 = ~pi13 & ~n2882;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = ~n2624 & n2756;
  assign n2887 = n2680 & ~n2790;
  assign n2888 = ~n2680 & n2790;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = ~n2756 & n2889;
  assign n2891 = ~n2886 & ~n2890;
  assign n2892 = pi12 & n2891;
  assign n2893 = ~pi12 & ~n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2609 & n2756;
  assign n2896 = n2682 & ~n2794;
  assign n2897 = ~n2682 & n2794;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = ~n2756 & n2898;
  assign n2900 = ~n2895 & ~n2899;
  assign n2901 = pi14 & n2900;
  assign n2902 = ~pi14 & ~n2900;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n2885 & n2894;
  assign n2905 = n2903 & n2904;
  assign n2906 = n2876 & n2905;
  assign n2907 = n2867 & n2906;
  assign n2908 = ~n2666 & n2756;
  assign n2909 = n2669 & ~n2786;
  assign n2910 = ~n2669 & n2786;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = ~n2756 & n2911;
  assign n2913 = ~n2908 & ~n2912;
  assign n2914 = pi10 & ~n2913;
  assign n2915 = ~pi10 & n2913;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = n2640 & n2756;
  assign n2918 = n2643 & ~n2788;
  assign n2919 = ~n2643 & n2788;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = ~n2756 & n2920;
  assign n2922 = ~n2917 & ~n2921;
  assign n2923 = pi11 & ~n2922;
  assign n2924 = ~pi11 & n2922;
  assign n2925 = ~n2923 & ~n2924;
  assign n2926 = ~pi08 & n2780;
  assign n2927 = ~n2649 & n2756;
  assign n2928 = n2652 & ~n2784;
  assign n2929 = ~n2652 & n2784;
  assign n2930 = ~n2928 & ~n2929;
  assign n2931 = ~n2756 & n2930;
  assign n2932 = ~n2927 & ~n2931;
  assign n2933 = pi09 & ~n2932;
  assign n2934 = ~pi09 & n2932;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n2916 & ~n2926;
  assign n2937 = n2925 & n2935;
  assign n2938 = n2936 & n2937;
  assign n2939 = ~n2781 & n2938;
  assign n2940 = n2907 & n2939;
  assign n2941 = n2697 & n2756;
  assign n2942 = n2743 & ~n2772;
  assign n2943 = ~n2743 & n2772;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n2756 & n2944;
  assign n2946 = ~n2941 & ~n2945;
  assign n2947 = pi07 & ~n2946;
  assign n2948 = ~n2705 & n2756;
  assign n2949 = n2744 & ~n2770;
  assign n2950 = ~n2744 & n2770;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = ~n2756 & n2951;
  assign n2953 = ~n2948 & ~n2952;
  assign n2954 = ~pi06 & n2953;
  assign n2955 = ~pi07 & n2946;
  assign n2956 = ~n2712 & n2756;
  assign n2957 = ~n2742 & ~n2768;
  assign n2958 = n2742 & n2768;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~n2756 & n2959;
  assign n2961 = ~n2956 & ~n2960;
  assign n2962 = pi05 & ~n2961;
  assign n2963 = pi06 & ~n2953;
  assign n2964 = ~pi05 & n2961;
  assign n2965 = n2721 & n2756;
  assign n2966 = n2746 & ~n2766;
  assign n2967 = ~n2746 & n2766;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = ~n2756 & n2968;
  assign n2970 = ~n2965 & ~n2969;
  assign n2971 = pi04 & ~n2970;
  assign n2972 = ~n2964 & n2971;
  assign n2973 = ~n2962 & ~n2963;
  assign n2974 = ~n2972 & n2973;
  assign n2975 = ~n2954 & ~n2955;
  assign n2976 = ~n2974 & n2975;
  assign n2977 = ~n2947 & ~n2976;
  assign n2978 = n2940 & n2977;
  assign n2979 = ~n2839 & ~n2848;
  assign n2980 = ~n2840 & ~n2979;
  assign n2981 = ~n2859 & n2980;
  assign n2982 = ~n2858 & ~n2981;
  assign n2983 = ~n2830 & n2982;
  assign n2984 = ~n2831 & ~n2983;
  assign n2985 = ~n2822 & n2984;
  assign n2986 = n74 & ~n2821;
  assign n2987 = ~n2985 & n2986;
  assign n2988 = ~n2866 & n2987;
  assign n2989 = ~n2884 & n2892;
  assign n2990 = ~n2883 & ~n2901;
  assign n2991 = ~n2989 & n2990;
  assign n2992 = ~n2875 & ~n2902;
  assign n2993 = ~n2991 & n2992;
  assign n2994 = ~n2874 & ~n2993;
  assign n2995 = n2867 & n2994;
  assign n2996 = ~n2907 & ~n2988;
  assign n2997 = ~n2995 & n2996;
  assign n2998 = ~n2914 & ~n2933;
  assign n2999 = ~n2915 & ~n2924;
  assign n3000 = ~n2998 & n2999;
  assign n3001 = ~n2923 & ~n3000;
  assign n3002 = ~n2938 & n3001;
  assign n3003 = n2907 & ~n3002;
  assign n3004 = ~n2997 & ~n3003;
  assign n3005 = ~n2978 & ~n3004;
  assign n3006 = ~n2954 & ~n2963;
  assign n3007 = ~n2962 & ~n2964;
  assign n3008 = ~n2947 & ~n2955;
  assign n3009 = ~pi04 & n2970;
  assign n3010 = ~n2971 & ~n3009;
  assign n3011 = n3006 & n3007;
  assign n3012 = n3008 & n3010;
  assign n3013 = n3011 & n3012;
  assign n3014 = n2940 & n3013;
  assign n3015 = n2736 & n2756;
  assign n3016 = ~n2753 & ~n2759;
  assign n3017 = n2753 & n2759;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~n2756 & n3018;
  assign n3020 = ~n3015 & ~n3019;
  assign n3021 = ~pi03 & ~n3020;
  assign n3022 = pi00 & ~n2756;
  assign n3023 = ~pi01 & n3022;
  assign n3024 = ~pi02 & n2763;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = pi02 & ~n2763;
  assign n3027 = pi03 & n3020;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = ~n3025 & n3028;
  assign n3030 = ~n3021 & ~n3029;
  assign n3031 = n3014 & n3030;
  assign n3032 = ~n3005 & ~n3031;
  assign n3033 = ~n3024 & ~n3026;
  assign n3034 = ~n3021 & ~n3027;
  assign n3035 = n84 & n3033;
  assign n3036 = n3034 & n3035;
  assign n3037 = n3014 & n3036;
  assign n3038 = ~n3032 & ~n3037;
  assign n3039 = ~n2763 & n3038;
  assign n3040 = ~n84 & ~n3023;
  assign n3041 = ~n3033 & ~n3040;
  assign n3042 = n3033 & n3040;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = ~n3038 & n3043;
  assign n3045 = ~n3039 & ~n3044;
  assign n3046 = pi03 & ~n3045;
  assign n3047 = ~pi03 & n3045;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = n3020 & n3038;
  assign n3050 = ~n3024 & n3040;
  assign n3051 = ~n3026 & ~n3050;
  assign n3052 = n3034 & ~n3051;
  assign n3053 = ~n3034 & n3051;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = ~n3038 & n3054;
  assign n3056 = ~n3049 & ~n3055;
  assign n3057 = pi04 & ~n3056;
  assign n3058 = ~pi04 & n3056;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = n2803 & n3038;
  assign n3061 = ~n2804 & ~n2851;
  assign n3062 = ~n3027 & n3051;
  assign n3063 = ~n3021 & ~n3062;
  assign n3064 = ~n3009 & n3063;
  assign n3065 = ~n2971 & ~n3064;
  assign n3066 = ~n2964 & ~n3065;
  assign n3067 = ~n2962 & ~n3066;
  assign n3068 = ~n2954 & ~n3067;
  assign n3069 = ~n2963 & ~n3068;
  assign n3070 = ~n2955 & ~n3069;
  assign n3071 = ~n2947 & ~n3070;
  assign n3072 = ~n2926 & ~n3071;
  assign n3073 = ~n2781 & ~n3072;
  assign n3074 = ~n2934 & ~n3073;
  assign n3075 = ~n2933 & ~n3074;
  assign n3076 = ~n2914 & n3075;
  assign n3077 = ~n2915 & ~n3076;
  assign n3078 = ~n2923 & ~n3077;
  assign n3079 = ~n2924 & ~n3078;
  assign n3080 = ~n2892 & ~n3079;
  assign n3081 = ~n2893 & ~n3080;
  assign n3082 = ~n2883 & ~n3081;
  assign n3083 = ~n2884 & ~n3082;
  assign n3084 = ~n2901 & ~n3083;
  assign n3085 = ~n2902 & ~n3084;
  assign n3086 = ~n2874 & ~n3085;
  assign n3087 = ~n2875 & ~n3086;
  assign n3088 = ~n3061 & ~n3087;
  assign n3089 = n3061 & n3087;
  assign n3090 = ~n3038 & ~n3088;
  assign n3091 = ~n3089 & n3090;
  assign n3092 = ~n3060 & ~n3091;
  assign n3093 = ~pi17 & n3092;
  assign n3094 = pi17 & ~n3092;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = ~n2820 & n3038;
  assign n3097 = ~n2804 & ~n3087;
  assign n3098 = ~n2851 & ~n3097;
  assign n3099 = ~n2849 & n3098;
  assign n3100 = ~n2848 & ~n3099;
  assign n3101 = ~n2839 & n3100;
  assign n3102 = ~n2840 & ~n3101;
  assign n3103 = ~n2859 & n3102;
  assign n3104 = ~n2858 & ~n3103;
  assign n3105 = ~n2831 & ~n3104;
  assign n3106 = ~n2830 & ~n3105;
  assign n3107 = n2823 & ~n3106;
  assign n3108 = ~n2823 & n3106;
  assign n3109 = ~n3038 & ~n3107;
  assign n3110 = ~n3108 & n3109;
  assign n3111 = ~n3096 & ~n3110;
  assign n3112 = pi22 & ~n3111;
  assign n3113 = ~pi22 & n3111;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = ~n2857 & n3038;
  assign n3116 = ~n2860 & ~n3102;
  assign n3117 = n2860 & n3102;
  assign n3118 = ~n3038 & ~n3116;
  assign n3119 = ~n3117 & n3118;
  assign n3120 = ~n3115 & ~n3119;
  assign n3121 = pi20 & ~n3120;
  assign n3122 = ~pi20 & n3120;
  assign n3123 = ~n3121 & ~n3122;
  assign n3124 = ~n2829 & n3038;
  assign n3125 = n2832 & ~n3104;
  assign n3126 = ~n2832 & n3104;
  assign n3127 = ~n3038 & ~n3125;
  assign n3128 = ~n3126 & n3127;
  assign n3129 = ~n3124 & ~n3128;
  assign n3130 = pi21 & ~n3129;
  assign n3131 = ~pi21 & n3129;
  assign n3132 = ~n3130 & ~n3131;
  assign n3133 = n2838 & n3038;
  assign n3134 = n2841 & ~n3100;
  assign n3135 = ~n2841 & n3100;
  assign n3136 = ~n3038 & ~n3134;
  assign n3137 = ~n3135 & n3136;
  assign n3138 = ~n3133 & ~n3137;
  assign n3139 = pi19 & ~n3138;
  assign n3140 = ~pi19 & n3138;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = ~n2847 & n3038;
  assign n3143 = ~n2850 & ~n3098;
  assign n3144 = n2850 & n3098;
  assign n3145 = ~n3038 & ~n3143;
  assign n3146 = ~n3144 & n3145;
  assign n3147 = ~n3142 & ~n3146;
  assign n3148 = pi18 & ~n3147;
  assign n3149 = ~pi18 & n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = n73 & n3150;
  assign n3152 = n3141 & n3151;
  assign n3153 = n3123 & n3152;
  assign n3154 = n3132 & n3153;
  assign n3155 = n3114 & n3154;
  assign n3156 = n3095 & n3155;
  assign n3157 = ~n2873 & n3038;
  assign n3158 = n2876 & ~n3085;
  assign n3159 = ~n2876 & n3085;
  assign n3160 = ~n3038 & ~n3158;
  assign n3161 = ~n3159 & n3160;
  assign n3162 = ~n3157 & ~n3161;
  assign n3163 = pi16 & n3162;
  assign n3164 = ~pi16 & ~n3162;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = ~n2882 & n3038;
  assign n3167 = n2885 & ~n3081;
  assign n3168 = ~n2885 & n3081;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~n3038 & n3169;
  assign n3171 = ~n3166 & ~n3170;
  assign n3172 = pi14 & n3171;
  assign n3173 = ~pi14 & ~n3171;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = ~n2891 & n3038;
  assign n3176 = n2894 & ~n3079;
  assign n3177 = ~n2894 & n3079;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~n3038 & n3178;
  assign n3180 = ~n3175 & ~n3179;
  assign n3181 = pi13 & n3180;
  assign n3182 = ~pi13 & ~n3180;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = ~n2900 & n3038;
  assign n3185 = n2903 & ~n3083;
  assign n3186 = ~n2903 & n3083;
  assign n3187 = ~n3038 & ~n3185;
  assign n3188 = ~n3186 & n3187;
  assign n3189 = ~n3184 & ~n3188;
  assign n3190 = ~pi15 & ~n3189;
  assign n3191 = pi15 & n3189;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = n3174 & n3183;
  assign n3194 = n3192 & n3193;
  assign n3195 = n3165 & n3194;
  assign n3196 = n3156 & n3195;
  assign n3197 = ~n2913 & n3038;
  assign n3198 = n2916 & ~n3075;
  assign n3199 = ~n2916 & n3075;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = ~n3038 & n3200;
  assign n3202 = ~n3197 & ~n3201;
  assign n3203 = ~pi11 & n3202;
  assign n3204 = pi11 & ~n3202;
  assign n3205 = ~n3203 & ~n3204;
  assign n3206 = ~n2932 & n3038;
  assign n3207 = n2935 & ~n3073;
  assign n3208 = ~n2935 & n3073;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = ~n3038 & n3209;
  assign n3211 = ~n3206 & ~n3210;
  assign n3212 = ~pi10 & n3211;
  assign n3213 = pi10 & ~n3211;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = ~n2781 & ~n2926;
  assign n3216 = ~n3071 & ~n3215;
  assign n3217 = n3071 & n3215;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = ~n3038 & ~n3218;
  assign n3220 = ~n2780 & n3038;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = ~pi09 & n3221;
  assign n3223 = pi09 & ~n3221;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = ~n2925 & ~n3077;
  assign n3226 = n2925 & n3077;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = ~n3038 & ~n3227;
  assign n3229 = n2922 & n3038;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = ~pi12 & ~n3230;
  assign n3232 = pi12 & n3230;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = n3205 & n3214;
  assign n3235 = n3224 & n3233;
  assign n3236 = n3234 & n3235;
  assign n3237 = n3196 & n3236;
  assign n3238 = ~n2946 & n3038;
  assign n3239 = n3008 & ~n3069;
  assign n3240 = ~n3008 & n3069;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~n3038 & n3241;
  assign n3243 = ~n3238 & ~n3242;
  assign n3244 = pi08 & ~n3243;
  assign n3245 = ~pi08 & n3243;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = ~n2953 & n3038;
  assign n3248 = n3006 & ~n3067;
  assign n3249 = ~n3006 & n3067;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = ~n3038 & n3250;
  assign n3252 = ~n3247 & ~n3251;
  assign n3253 = pi07 & ~n3252;
  assign n3254 = ~pi07 & n3252;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = ~n3007 & ~n3065;
  assign n3257 = n3007 & n3065;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = ~n3038 & ~n3258;
  assign n3260 = ~n2961 & n3038;
  assign n3261 = ~n3259 & ~n3260;
  assign n3262 = pi06 & ~n3261;
  assign n3263 = ~pi06 & n3261;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = n2970 & n3038;
  assign n3266 = n3010 & ~n3063;
  assign n3267 = ~n3010 & n3063;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = ~n3038 & n3268;
  assign n3270 = ~n3265 & ~n3269;
  assign n3271 = pi05 & n3270;
  assign n3272 = ~pi05 & ~n3270;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = n3246 & n3255;
  assign n3275 = n3264 & n3273;
  assign n3276 = n3274 & n3275;
  assign n3277 = n3237 & n3276;
  assign n3278 = n3048 & n3059;
  assign n3279 = n3277 & n3278;
  assign n3280 = pi00 & ~n2752;
  assign n3281 = ~pi01 & ~n3280;
  assign n3282 = pi01 & n3280;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = ~n3038 & ~n3283;
  assign n3285 = ~n3022 & n3038;
  assign n3286 = ~n3284 & ~n3285;
  assign n3287 = pi02 & ~n3286;
  assign n3288 = ~pi02 & n3286;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = pi00 & ~n3038;
  assign n3291 = ~pi01 & n3290;
  assign n3292 = n3289 & ~n3291;
  assign n3293 = n3279 & n3292;
  assign n3294 = ~n3172 & ~n3181;
  assign n3295 = ~n3173 & ~n3294;
  assign n3296 = ~n3190 & n3295;
  assign n3297 = ~n3191 & ~n3296;
  assign n3298 = ~n3163 & n3297;
  assign n3299 = ~n3164 & ~n3298;
  assign n3300 = n3156 & ~n3299;
  assign n3301 = ~n3093 & n3155;
  assign n3302 = ~n3139 & ~n3148;
  assign n3303 = ~n3140 & ~n3302;
  assign n3304 = ~n3122 & n3303;
  assign n3305 = ~n3121 & ~n3304;
  assign n3306 = ~n3130 & n3305;
  assign n3307 = ~n3131 & ~n3306;
  assign n3308 = ~n3113 & n3307;
  assign n3309 = n73 & ~n3112;
  assign n3310 = ~n3308 & n3309;
  assign n3311 = ~n3301 & n3310;
  assign n3312 = ~n3300 & ~n3311;
  assign n3313 = ~n3213 & n3222;
  assign n3314 = ~n3203 & ~n3212;
  assign n3315 = ~n3313 & n3314;
  assign n3316 = ~n3204 & ~n3315;
  assign n3317 = ~n3231 & ~n3316;
  assign n3318 = ~n3232 & ~n3317;
  assign n3319 = n3196 & ~n3318;
  assign n3320 = ~n3312 & ~n3319;
  assign n3321 = ~n3262 & ~n3271;
  assign n3322 = ~n3254 & ~n3263;
  assign n3323 = ~n3321 & n3322;
  assign n3324 = ~n3244 & ~n3253;
  assign n3325 = ~n3323 & n3324;
  assign n3326 = ~n3245 & ~n3325;
  assign n3327 = n3237 & ~n3326;
  assign n3328 = ~n3320 & ~n3327;
  assign n3329 = ~n3047 & n3287;
  assign n3330 = ~n3046 & ~n3057;
  assign n3331 = ~n3329 & n3330;
  assign n3332 = ~n3058 & ~n3331;
  assign n3333 = n3277 & n3332;
  assign n3334 = ~n3328 & ~n3333;
  assign n3335 = ~n3293 & n3334;
  assign n3336 = n84 & n3289;
  assign n3337 = n3279 & n3336;
  assign n3338 = ~n3335 & ~n3337;
  assign n3339 = pi01 & n3032;
  assign n3340 = n314 & ~n3032;
  assign n3341 = ~n3339 & ~n3340;
  assign n3342 = ~n3338 & n3341;
  assign n3343 = ~n3290 & n3338;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = ~pi02 & n3344;
  assign n3346 = n3180 & n3338;
  assign n3347 = ~n84 & ~n3291;
  assign n3348 = ~n3287 & ~n3347;
  assign n3349 = ~n3288 & ~n3348;
  assign n3350 = ~n3047 & n3349;
  assign n3351 = ~n3046 & ~n3350;
  assign n3352 = ~n3057 & n3351;
  assign n3353 = ~n3058 & ~n3352;
  assign n3354 = ~n3271 & ~n3353;
  assign n3355 = ~n3272 & ~n3354;
  assign n3356 = ~n3262 & ~n3355;
  assign n3357 = ~n3263 & ~n3356;
  assign n3358 = ~n3254 & n3357;
  assign n3359 = ~n3253 & ~n3358;
  assign n3360 = ~n3245 & ~n3359;
  assign n3361 = ~n3244 & ~n3360;
  assign n3362 = ~n3222 & ~n3361;
  assign n3363 = ~n3223 & ~n3362;
  assign n3364 = ~n3212 & ~n3363;
  assign n3365 = ~n3213 & ~n3364;
  assign n3366 = ~n3203 & ~n3365;
  assign n3367 = ~n3204 & ~n3366;
  assign n3368 = ~n3231 & ~n3367;
  assign n3369 = ~n3232 & ~n3368;
  assign n3370 = n3183 & ~n3369;
  assign n3371 = ~n3183 & n3369;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = ~n3338 & n3372;
  assign n3374 = ~n3346 & ~n3373;
  assign n3375 = pi14 & ~n3374;
  assign n3376 = ~pi14 & n3374;
  assign n3377 = ~n3375 & ~n3376;
  assign n3378 = ~n3181 & n3369;
  assign n3379 = ~n3182 & ~n3378;
  assign n3380 = ~n3174 & ~n3379;
  assign n3381 = n3174 & n3379;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = ~n3338 & ~n3382;
  assign n3384 = ~n3171 & n3338;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = pi15 & n3385;
  assign n3387 = ~pi15 & ~n3385;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = ~n3172 & ~n3379;
  assign n3390 = ~n3173 & ~n3389;
  assign n3391 = ~n3191 & ~n3390;
  assign n3392 = ~n3190 & ~n3391;
  assign n3393 = ~n3165 & ~n3392;
  assign n3394 = n3165 & n3392;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = ~n3338 & ~n3395;
  assign n3397 = ~n3162 & n3338;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = pi17 & n3398;
  assign n3400 = ~pi17 & ~n3398;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = n3092 & n3338;
  assign n3403 = ~n3163 & ~n3392;
  assign n3404 = ~n3164 & ~n3403;
  assign n3405 = n3095 & ~n3404;
  assign n3406 = ~n3095 & n3404;
  assign n3407 = ~n3338 & ~n3405;
  assign n3408 = ~n3406 & n3407;
  assign n3409 = ~n3402 & ~n3408;
  assign n3410 = pi18 & n3409;
  assign n3411 = n3147 & n3338;
  assign n3412 = ~n3094 & ~n3404;
  assign n3413 = ~n3093 & ~n3412;
  assign n3414 = n3150 & ~n3413;
  assign n3415 = ~n3150 & n3413;
  assign n3416 = ~n3338 & ~n3414;
  assign n3417 = ~n3415 & n3416;
  assign n3418 = ~n3411 & ~n3417;
  assign n3419 = pi19 & n3418;
  assign n3420 = ~pi19 & ~n3418;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = ~n3120 & n3338;
  assign n3423 = ~n3148 & ~n3413;
  assign n3424 = ~n3149 & ~n3423;
  assign n3425 = ~n3140 & n3424;
  assign n3426 = ~n3139 & ~n3425;
  assign n3427 = n3123 & ~n3426;
  assign n3428 = ~n3123 & n3426;
  assign n3429 = ~n3338 & ~n3427;
  assign n3430 = ~n3428 & n3429;
  assign n3431 = ~n3422 & ~n3430;
  assign n3432 = pi21 & ~n3431;
  assign n3433 = ~pi21 & n3431;
  assign n3434 = ~n3432 & ~n3433;
  assign n3435 = ~pi18 & ~n3409;
  assign n3436 = ~pi24 & n71;
  assign n3437 = ~n3138 & n3338;
  assign n3438 = ~n3141 & ~n3424;
  assign n3439 = n3141 & n3424;
  assign n3440 = ~n3338 & ~n3438;
  assign n3441 = ~n3439 & n3440;
  assign n3442 = ~n3437 & ~n3441;
  assign n3443 = pi20 & ~n3442;
  assign n3444 = ~pi20 & n3442;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = ~n3111 & n3338;
  assign n3447 = ~n3122 & ~n3426;
  assign n3448 = ~n3121 & ~n3447;
  assign n3449 = ~n3131 & ~n3448;
  assign n3450 = ~n3130 & ~n3449;
  assign n3451 = n3114 & ~n3450;
  assign n3452 = ~n3114 & n3450;
  assign n3453 = ~n3338 & ~n3451;
  assign n3454 = ~n3452 & n3453;
  assign n3455 = ~n3446 & ~n3454;
  assign n3456 = pi23 & ~n3455;
  assign n3457 = ~pi23 & n3455;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = ~n3129 & n3338;
  assign n3460 = n3132 & ~n3448;
  assign n3461 = ~n3132 & n3448;
  assign n3462 = ~n3338 & ~n3460;
  assign n3463 = ~n3461 & n3462;
  assign n3464 = ~n3459 & ~n3463;
  assign n3465 = pi22 & ~n3464;
  assign n3466 = ~pi22 & n3464;
  assign n3467 = ~n3465 & ~n3466;
  assign n3468 = ~n3435 & n3436;
  assign n3469 = n3421 & n3468;
  assign n3470 = n3445 & n3469;
  assign n3471 = n3434 & n3470;
  assign n3472 = n3467 & n3471;
  assign n3473 = n3458 & n3472;
  assign n3474 = ~n3410 & n3473;
  assign n3475 = ~n3192 & ~n3390;
  assign n3476 = n3192 & n3390;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = ~n3338 & ~n3477;
  assign n3479 = ~n3189 & n3338;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = pi16 & n3480;
  assign n3482 = ~pi16 & ~n3480;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = n3377 & n3388;
  assign n3485 = n3483 & n3484;
  assign n3486 = n3401 & n3485;
  assign n3487 = n3474 & n3486;
  assign n3488 = ~n3211 & n3338;
  assign n3489 = n3214 & ~n3363;
  assign n3490 = ~n3214 & n3363;
  assign n3491 = ~n3489 & ~n3490;
  assign n3492 = ~n3338 & n3491;
  assign n3493 = ~n3488 & ~n3492;
  assign n3494 = ~pi11 & n3493;
  assign n3495 = pi11 & ~n3493;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = ~n3202 & n3338;
  assign n3498 = n3205 & ~n3365;
  assign n3499 = ~n3205 & n3365;
  assign n3500 = ~n3498 & ~n3499;
  assign n3501 = ~n3338 & n3500;
  assign n3502 = ~n3497 & ~n3501;
  assign n3503 = ~pi12 & n3502;
  assign n3504 = pi12 & ~n3502;
  assign n3505 = ~n3503 & ~n3504;
  assign n3506 = ~n3233 & ~n3367;
  assign n3507 = n3233 & n3367;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~n3338 & ~n3508;
  assign n3510 = n3230 & n3338;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = pi13 & ~n3511;
  assign n3513 = ~pi13 & n3511;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = ~n3221 & n3338;
  assign n3516 = n3224 & ~n3361;
  assign n3517 = ~n3224 & n3361;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = ~n3338 & n3518;
  assign n3520 = ~n3515 & ~n3519;
  assign n3521 = ~pi10 & n3520;
  assign n3522 = pi10 & ~n3520;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = n3496 & n3505;
  assign n3525 = n3514 & n3523;
  assign n3526 = n3524 & n3525;
  assign n3527 = n3487 & n3526;
  assign n3528 = n3261 & n3338;
  assign n3529 = n3264 & ~n3355;
  assign n3530 = ~n3264 & n3355;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~n3338 & n3531;
  assign n3533 = ~n3528 & ~n3532;
  assign n3534 = pi07 & n3533;
  assign n3535 = ~pi07 & ~n3533;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = ~n3243 & n3338;
  assign n3538 = n3246 & ~n3359;
  assign n3539 = ~n3246 & n3359;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = ~n3338 & n3540;
  assign n3542 = ~n3537 & ~n3541;
  assign n3543 = pi09 & ~n3542;
  assign n3544 = ~pi09 & n3542;
  assign n3545 = ~n3543 & ~n3544;
  assign n3546 = n3252 & n3338;
  assign n3547 = n3255 & ~n3357;
  assign n3548 = ~n3255 & n3357;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = ~n3338 & n3549;
  assign n3551 = ~n3546 & ~n3550;
  assign n3552 = pi08 & n3551;
  assign n3553 = ~pi08 & ~n3551;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = ~n3273 & ~n3353;
  assign n3556 = n3273 & n3353;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = ~n3338 & ~n3557;
  assign n3559 = ~n3270 & n3338;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = pi06 & n3560;
  assign n3562 = ~pi06 & ~n3560;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = n3536 & n3545;
  assign n3565 = n3554 & n3563;
  assign n3566 = n3564 & n3565;
  assign n3567 = n3527 & n3566;
  assign n3568 = ~n3045 & n3338;
  assign n3569 = ~n3048 & ~n3349;
  assign n3570 = n3048 & n3349;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3338 & n3571;
  assign n3573 = ~n3568 & ~n3572;
  assign n3574 = ~pi04 & n3573;
  assign n3575 = pi04 & ~n3573;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~n3286 & n3338;
  assign n3578 = ~n3289 & ~n3347;
  assign n3579 = n3289 & n3347;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = ~n3338 & n3580;
  assign n3582 = ~n3577 & ~n3581;
  assign n3583 = pi03 & ~n3582;
  assign n3584 = ~pi03 & n3582;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = ~n3056 & n3338;
  assign n3587 = n3059 & ~n3351;
  assign n3588 = ~n3059 & n3351;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3338 & n3589;
  assign n3591 = ~n3586 & ~n3590;
  assign n3592 = ~pi05 & n3591;
  assign n3593 = pi05 & ~n3591;
  assign n3594 = ~n3592 & ~n3593;
  assign n3595 = n3576 & n3585;
  assign n3596 = n3594 & n3595;
  assign n3597 = n3567 & n3596;
  assign n3598 = ~n3345 & n3597;
  assign n3599 = ~n3494 & ~n3521;
  assign n3600 = ~n3495 & ~n3504;
  assign n3601 = ~n3599 & n3600;
  assign n3602 = ~n3503 & ~n3513;
  assign n3603 = ~n3601 & n3602;
  assign n3604 = ~n3512 & ~n3603;
  assign n3605 = n3487 & ~n3604;
  assign n3606 = ~n3419 & ~n3443;
  assign n3607 = ~n3444 & ~n3606;
  assign n3608 = ~n3432 & ~n3607;
  assign n3609 = ~n3433 & ~n3608;
  assign n3610 = ~n3465 & ~n3609;
  assign n3611 = ~n3466 & ~n3610;
  assign n3612 = ~n3457 & n3611;
  assign n3613 = n3436 & ~n3456;
  assign n3614 = ~n3612 & n3613;
  assign n3615 = ~n3473 & n3614;
  assign n3616 = n3375 & ~n3387;
  assign n3617 = ~n3386 & ~n3616;
  assign n3618 = ~n3481 & n3617;
  assign n3619 = ~n3482 & ~n3618;
  assign n3620 = ~n3400 & n3619;
  assign n3621 = ~n3399 & ~n3620;
  assign n3622 = n3474 & n3621;
  assign n3623 = ~n3615 & ~n3622;
  assign n3624 = ~n3605 & ~n3623;
  assign n3625 = ~n3534 & ~n3561;
  assign n3626 = ~n3535 & ~n3553;
  assign n3627 = ~n3625 & n3626;
  assign n3628 = ~n3543 & ~n3552;
  assign n3629 = ~n3627 & n3628;
  assign n3630 = ~n3544 & ~n3629;
  assign n3631 = n3527 & ~n3630;
  assign n3632 = ~n3624 & ~n3631;
  assign n3633 = ~n3575 & ~n3583;
  assign n3634 = ~n3574 & ~n3592;
  assign n3635 = ~n3633 & n3634;
  assign n3636 = ~n3593 & ~n3635;
  assign n3637 = n3567 & ~n3636;
  assign n3638 = ~n3632 & ~n3637;
  assign n3639 = ~n3598 & n3638;
  assign n3640 = pi02 & ~n3344;
  assign n3641 = ~n3345 & ~n3640;
  assign n3642 = n3597 & n3641;
  assign n3643 = pi00 & n3338;
  assign n3644 = ~pi01 & ~n3643;
  assign n3645 = n3642 & n3644;
  assign n3646 = ~n3639 & ~n3645;
  assign n3647 = pi00 & ~n3335;
  assign n3648 = ~pi01 & ~n3647;
  assign n3649 = pi01 & n3647;
  assign n3650 = ~n3648 & ~n3649;
  assign n3651 = ~n3646 & ~n3650;
  assign n3652 = pi00 & ~n3338;
  assign n3653 = n3646 & ~n3652;
  assign n3654 = ~n3651 & ~n3653;
  assign n3655 = n3542 & n3646;
  assign n3656 = ~n3345 & ~n3644;
  assign n3657 = ~n3640 & ~n3656;
  assign n3658 = ~n3584 & ~n3657;
  assign n3659 = ~n3583 & ~n3658;
  assign n3660 = ~n3575 & n3659;
  assign n3661 = ~n3574 & ~n3660;
  assign n3662 = ~n3592 & n3661;
  assign n3663 = ~n3593 & ~n3662;
  assign n3664 = ~n3561 & n3663;
  assign n3665 = ~n3562 & ~n3664;
  assign n3666 = ~n3534 & ~n3665;
  assign n3667 = ~n3535 & ~n3666;
  assign n3668 = ~n3552 & ~n3667;
  assign n3669 = ~n3553 & ~n3668;
  assign n3670 = n3545 & ~n3669;
  assign n3671 = ~n3545 & n3669;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = ~n3646 & n3672;
  assign n3674 = ~n3655 & ~n3673;
  assign n3675 = pi10 & n3674;
  assign n3676 = ~pi10 & ~n3674;
  assign n3677 = ~n3551 & n3646;
  assign n3678 = n3554 & ~n3667;
  assign n3679 = ~n3554 & n3667;
  assign n3680 = ~n3678 & ~n3679;
  assign n3681 = ~n3646 & n3680;
  assign n3682 = ~n3677 & ~n3681;
  assign n3683 = pi09 & n3682;
  assign n3684 = ~n3533 & n3646;
  assign n3685 = n3536 & ~n3665;
  assign n3686 = ~n3536 & n3665;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = ~n3646 & n3687;
  assign n3689 = ~n3684 & ~n3688;
  assign n3690 = pi08 & n3689;
  assign n3691 = ~n3563 & ~n3663;
  assign n3692 = n3563 & n3663;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = ~n3646 & ~n3693;
  assign n3695 = n3560 & n3646;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = pi07 & ~n3696;
  assign n3698 = ~n3690 & ~n3697;
  assign n3699 = ~pi08 & ~n3689;
  assign n3700 = ~pi09 & ~n3682;
  assign n3701 = ~n3699 & ~n3700;
  assign n3702 = ~n3698 & n3701;
  assign n3703 = ~n3683 & ~n3702;
  assign n3704 = ~n3676 & ~n3703;
  assign n3705 = n3409 & n3646;
  assign n3706 = ~n3543 & ~n3669;
  assign n3707 = ~n3544 & ~n3706;
  assign n3708 = ~n3522 & ~n3707;
  assign n3709 = n3599 & ~n3708;
  assign n3710 = n3600 & ~n3709;
  assign n3711 = ~n3503 & ~n3710;
  assign n3712 = ~n3513 & n3711;
  assign n3713 = ~n3512 & ~n3712;
  assign n3714 = ~n3376 & ~n3713;
  assign n3715 = ~n3375 & ~n3714;
  assign n3716 = ~n3387 & ~n3715;
  assign n3717 = ~n3386 & ~n3716;
  assign n3718 = ~n3481 & n3717;
  assign n3719 = ~n3482 & ~n3718;
  assign n3720 = ~n3399 & ~n3719;
  assign n3721 = ~n3400 & ~n3720;
  assign n3722 = ~n3410 & ~n3435;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = n3721 & n3722;
  assign n3725 = ~n3646 & ~n3723;
  assign n3726 = ~n3724 & n3725;
  assign n3727 = ~n3705 & ~n3726;
  assign n3728 = pi19 & ~n3727;
  assign n3729 = ~pi19 & n3727;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = ~n3455 & n3646;
  assign n3732 = ~n3410 & ~n3721;
  assign n3733 = ~n3435 & ~n3732;
  assign n3734 = ~n3419 & ~n3733;
  assign n3735 = ~n3420 & ~n3734;
  assign n3736 = ~n3444 & n3735;
  assign n3737 = ~n3443 & ~n3736;
  assign n3738 = ~n3433 & ~n3737;
  assign n3739 = ~n3432 & ~n3738;
  assign n3740 = ~n3466 & ~n3739;
  assign n3741 = ~n3465 & ~n3740;
  assign n3742 = n3458 & ~n3741;
  assign n3743 = ~n3458 & n3741;
  assign n3744 = ~n3646 & ~n3742;
  assign n3745 = ~n3743 & n3744;
  assign n3746 = ~n3731 & ~n3745;
  assign n3747 = pi24 & ~n3746;
  assign n3748 = ~pi24 & n3746;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = ~n3431 & n3646;
  assign n3751 = n3434 & ~n3737;
  assign n3752 = ~n3434 & n3737;
  assign n3753 = ~n3646 & ~n3751;
  assign n3754 = ~n3752 & n3753;
  assign n3755 = ~n3750 & ~n3754;
  assign n3756 = pi22 & ~n3755;
  assign n3757 = ~pi22 & n3755;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = ~n3464 & n3646;
  assign n3760 = n3467 & ~n3739;
  assign n3761 = ~n3467 & n3739;
  assign n3762 = ~n3646 & ~n3760;
  assign n3763 = ~n3761 & n3762;
  assign n3764 = ~n3759 & ~n3763;
  assign n3765 = pi23 & ~n3764;
  assign n3766 = ~pi23 & n3764;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = n3442 & n3646;
  assign n3769 = n3445 & ~n3735;
  assign n3770 = ~n3445 & n3735;
  assign n3771 = ~n3646 & ~n3769;
  assign n3772 = ~n3770 & n3771;
  assign n3773 = ~n3768 & ~n3772;
  assign n3774 = pi21 & n3773;
  assign n3775 = ~pi21 & ~n3773;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = ~n3421 & ~n3733;
  assign n3778 = n3421 & n3733;
  assign n3779 = ~n3777 & ~n3778;
  assign n3780 = ~n3646 & ~n3779;
  assign n3781 = ~n3418 & n3646;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = pi20 & n3782;
  assign n3784 = ~pi20 & ~n3782;
  assign n3785 = ~n3783 & ~n3784;
  assign n3786 = n71 & n3785;
  assign n3787 = n3776 & n3786;
  assign n3788 = n3758 & n3787;
  assign n3789 = n3767 & n3788;
  assign n3790 = n3749 & n3789;
  assign n3791 = n3730 & n3790;
  assign n3792 = ~n3401 & ~n3719;
  assign n3793 = n3401 & n3719;
  assign n3794 = ~n3792 & ~n3793;
  assign n3795 = ~n3646 & ~n3794;
  assign n3796 = ~n3398 & n3646;
  assign n3797 = ~n3795 & ~n3796;
  assign n3798 = pi18 & n3797;
  assign n3799 = ~pi18 & ~n3797;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = ~n3374 & n3646;
  assign n3802 = n3377 & ~n3713;
  assign n3803 = ~n3377 & n3713;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = ~n3646 & n3804;
  assign n3806 = ~n3801 & ~n3805;
  assign n3807 = pi15 & ~n3806;
  assign n3808 = ~pi15 & n3806;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = n3385 & n3646;
  assign n3811 = n3388 & ~n3715;
  assign n3812 = ~n3388 & n3715;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = ~n3646 & n3813;
  assign n3815 = ~n3810 & ~n3814;
  assign n3816 = pi16 & ~n3815;
  assign n3817 = ~pi16 & n3815;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = n3480 & n3646;
  assign n3820 = n3483 & ~n3717;
  assign n3821 = ~n3483 & n3717;
  assign n3822 = ~n3646 & ~n3820;
  assign n3823 = ~n3821 & n3822;
  assign n3824 = ~n3819 & ~n3823;
  assign n3825 = pi17 & ~n3824;
  assign n3826 = ~pi17 & n3824;
  assign n3827 = ~n3825 & ~n3826;
  assign n3828 = n3809 & n3818;
  assign n3829 = n3827 & n3828;
  assign n3830 = n3800 & n3829;
  assign n3831 = n3791 & n3830;
  assign n3832 = ~n3521 & ~n3708;
  assign n3833 = n3496 & ~n3832;
  assign n3834 = ~n3496 & n3832;
  assign n3835 = ~n3833 & ~n3834;
  assign n3836 = ~n3646 & ~n3835;
  assign n3837 = ~n3493 & n3646;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = pi12 & ~n3838;
  assign n3840 = ~pi12 & n3838;
  assign n3841 = ~n3839 & ~n3840;
  assign n3842 = n3520 & n3646;
  assign n3843 = n3523 & ~n3707;
  assign n3844 = ~n3523 & n3707;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = ~n3646 & n3845;
  assign n3847 = ~n3842 & ~n3846;
  assign n3848 = pi11 & n3847;
  assign n3849 = ~pi11 & ~n3847;
  assign n3850 = ~n3848 & ~n3849;
  assign n3851 = ~n3502 & n3646;
  assign n3852 = ~n3495 & ~n3709;
  assign n3853 = n3505 & ~n3852;
  assign n3854 = ~n3505 & n3852;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = ~n3646 & n3855;
  assign n3857 = ~n3851 & ~n3856;
  assign n3858 = pi13 & ~n3857;
  assign n3859 = ~pi13 & n3857;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = ~n3511 & n3646;
  assign n3862 = ~n3514 & ~n3711;
  assign n3863 = n3514 & n3711;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = ~n3646 & n3864;
  assign n3866 = ~n3861 & ~n3865;
  assign n3867 = pi14 & ~n3866;
  assign n3868 = ~pi14 & n3866;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = n3841 & n3850;
  assign n3871 = n3860 & n3869;
  assign n3872 = n3870 & n3871;
  assign n3873 = n3831 & n3872;
  assign n3874 = ~n3675 & ~n3704;
  assign n3875 = n3873 & n3874;
  assign n3876 = n3807 & ~n3817;
  assign n3877 = ~n3816 & ~n3876;
  assign n3878 = ~n3825 & n3877;
  assign n3879 = ~n3826 & ~n3878;
  assign n3880 = ~n3799 & n3879;
  assign n3881 = ~n3798 & ~n3880;
  assign n3882 = n3791 & n3881;
  assign n3883 = ~n3729 & n3790;
  assign n3884 = ~n3774 & ~n3783;
  assign n3885 = ~n3775 & ~n3884;
  assign n3886 = ~n3757 & n3885;
  assign n3887 = ~n3756 & ~n3886;
  assign n3888 = ~n3765 & n3887;
  assign n3889 = ~n3766 & ~n3888;
  assign n3890 = ~n3748 & n3889;
  assign n3891 = n71 & ~n3747;
  assign n3892 = ~n3890 & n3891;
  assign n3893 = ~n3883 & n3892;
  assign n3894 = ~n3882 & ~n3893;
  assign n3895 = ~n3840 & ~n3849;
  assign n3896 = ~n3839 & ~n3858;
  assign n3897 = ~n3895 & n3896;
  assign n3898 = ~n3859 & ~n3868;
  assign n3899 = ~n3897 & n3898;
  assign n3900 = ~n3867 & ~n3899;
  assign n3901 = n3831 & ~n3900;
  assign n3902 = ~n3894 & ~n3901;
  assign n3903 = ~n3875 & ~n3902;
  assign n3904 = ~n3591 & n3646;
  assign n3905 = ~n3594 & ~n3661;
  assign n3906 = n3594 & n3661;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = ~n3646 & n3907;
  assign n3909 = ~n3904 & ~n3908;
  assign n3910 = ~pi06 & n3909;
  assign n3911 = pi06 & ~n3909;
  assign n3912 = ~n3573 & n3646;
  assign n3913 = n3576 & ~n3659;
  assign n3914 = ~n3576 & n3659;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = ~n3646 & n3915;
  assign n3917 = ~n3912 & ~n3916;
  assign n3918 = ~pi05 & n3917;
  assign n3919 = ~n3582 & n3646;
  assign n3920 = n3585 & ~n3657;
  assign n3921 = ~n3585 & n3657;
  assign n3922 = ~n3920 & ~n3921;
  assign n3923 = ~n3646 & n3922;
  assign n3924 = ~n3919 & ~n3923;
  assign n3925 = ~pi04 & n3924;
  assign n3926 = n3344 & n3646;
  assign n3927 = ~n3641 & ~n3644;
  assign n3928 = n3641 & n3644;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~n3646 & n3929;
  assign n3931 = ~n3926 & ~n3930;
  assign n3932 = pi03 & n3931;
  assign n3933 = ~n3925 & n3932;
  assign n3934 = pi04 & ~n3924;
  assign n3935 = pi05 & ~n3917;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = ~n3933 & n3936;
  assign n3938 = ~n3918 & ~n3937;
  assign n3939 = ~n3911 & ~n3938;
  assign n3940 = ~n3675 & ~n3676;
  assign n3941 = ~n3683 & ~n3700;
  assign n3942 = ~n3690 & ~n3699;
  assign n3943 = ~pi07 & n3696;
  assign n3944 = ~n3697 & ~n3943;
  assign n3945 = n3940 & n3941;
  assign n3946 = n3942 & n3944;
  assign n3947 = n3945 & n3946;
  assign n3948 = n3873 & n3947;
  assign n3949 = ~n3910 & ~n3939;
  assign n3950 = n3948 & n3949;
  assign n3951 = ~n3903 & ~n3950;
  assign n3952 = ~n3910 & ~n3911;
  assign n3953 = ~n3925 & ~n3934;
  assign n3954 = ~pi03 & ~n3931;
  assign n3955 = ~n3932 & ~n3954;
  assign n3956 = ~n3918 & ~n3935;
  assign n3957 = n3952 & n3953;
  assign n3958 = n3955 & n3956;
  assign n3959 = n3957 & n3958;
  assign n3960 = n3948 & n3959;
  assign n3961 = ~n3951 & ~n3960;
  assign n3962 = pi02 & ~n3654;
  assign n3963 = ~pi02 & n3654;
  assign n3964 = pi00 & ~n3646;
  assign n3965 = ~pi01 & n3964;
  assign n3966 = ~n3963 & ~n3965;
  assign n3967 = ~n3962 & ~n3966;
  assign n3968 = n3960 & ~n3967;
  assign n3969 = ~n3961 & ~n3968;
  assign n3970 = ~n3962 & ~n3963;
  assign n3971 = n84 & n3970;
  assign n3972 = n3960 & n3971;
  assign n3973 = ~n3969 & ~n3972;
  assign n3974 = ~n3654 & n3973;
  assign n3975 = ~n84 & ~n3965;
  assign n3976 = ~n3970 & ~n3975;
  assign n3977 = n3970 & n3975;
  assign n3978 = ~n3976 & ~n3977;
  assign n3979 = ~n3973 & n3978;
  assign n3980 = ~n3974 & ~n3979;
  assign n3981 = ~n3917 & n3973;
  assign n3982 = ~n3962 & ~n3975;
  assign n3983 = ~n3963 & ~n3982;
  assign n3984 = ~n3932 & ~n3983;
  assign n3985 = ~n3954 & ~n3984;
  assign n3986 = ~n3925 & n3985;
  assign n3987 = ~n3934 & ~n3986;
  assign n3988 = n3956 & ~n3987;
  assign n3989 = ~n3956 & n3987;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = ~n3973 & n3990;
  assign n3992 = ~n3981 & ~n3991;
  assign n3993 = pi06 & ~n3992;
  assign n3994 = ~pi06 & n3992;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3764 & n3973;
  assign n3997 = ~n3935 & n3987;
  assign n3998 = ~n3918 & ~n3997;
  assign n3999 = ~n3910 & n3998;
  assign n4000 = ~n3911 & ~n3999;
  assign n4001 = ~n3943 & ~n4000;
  assign n4002 = ~n3697 & ~n4001;
  assign n4003 = ~n3690 & n4002;
  assign n4004 = ~n3699 & ~n4003;
  assign n4005 = ~n3683 & ~n4004;
  assign n4006 = ~n3700 & ~n4005;
  assign n4007 = ~n3675 & ~n4006;
  assign n4008 = ~n3676 & ~n4007;
  assign n4009 = ~n3848 & ~n4008;
  assign n4010 = ~n3849 & ~n4009;
  assign n4011 = ~n3840 & n4010;
  assign n4012 = ~n3839 & ~n4011;
  assign n4013 = ~n3859 & ~n4012;
  assign n4014 = ~n3858 & ~n4013;
  assign n4015 = ~n3868 & ~n4014;
  assign n4016 = ~n3867 & ~n4015;
  assign n4017 = ~n3808 & ~n4016;
  assign n4018 = ~n3807 & ~n4017;
  assign n4019 = ~n3817 & ~n4018;
  assign n4020 = ~n3816 & ~n4019;
  assign n4021 = ~n3825 & n4020;
  assign n4022 = ~n3826 & ~n4021;
  assign n4023 = ~n3798 & ~n4022;
  assign n4024 = ~n3799 & ~n4023;
  assign n4025 = ~n3728 & ~n4024;
  assign n4026 = ~n3729 & ~n4025;
  assign n4027 = ~n3783 & ~n4026;
  assign n4028 = ~n3784 & ~n4027;
  assign n4029 = ~n3774 & ~n4028;
  assign n4030 = ~n3775 & ~n4029;
  assign n4031 = ~n3756 & ~n4030;
  assign n4032 = ~n3757 & ~n4031;
  assign n4033 = ~n3767 & ~n4032;
  assign n4034 = n3767 & n4032;
  assign n4035 = ~n3973 & ~n4033;
  assign n4036 = ~n4034 & n4035;
  assign n4037 = ~n3996 & ~n4036;
  assign n4038 = pi24 & ~n4037;
  assign n4039 = ~pi24 & n4037;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = ~n3758 & ~n4030;
  assign n4042 = n3758 & n4030;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = ~n3973 & ~n4043;
  assign n4045 = n3755 & n3973;
  assign n4046 = ~n4044 & ~n4045;
  assign n4047 = pi23 & n4046;
  assign n4048 = ~pi23 & ~n4046;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = ~n3746 & n3973;
  assign n4051 = ~n3766 & n4032;
  assign n4052 = ~n3765 & ~n4051;
  assign n4053 = n3749 & ~n4052;
  assign n4054 = ~n3749 & n4052;
  assign n4055 = ~n3973 & ~n4053;
  assign n4056 = ~n4054 & n4055;
  assign n4057 = ~n4050 & ~n4056;
  assign n4058 = pi25 & ~n4057;
  assign n4059 = ~pi25 & n4057;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = ~n3773 & n3973;
  assign n4062 = n3776 & ~n4028;
  assign n4063 = ~n3776 & n4028;
  assign n4064 = ~n3973 & ~n4062;
  assign n4065 = ~n4063 & n4064;
  assign n4066 = ~n4061 & ~n4065;
  assign n4067 = pi22 & n4066;
  assign n4068 = ~pi22 & ~n4066;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = ~pi28 & n67;
  assign n4071 = ~pi27 & n4070;
  assign n4072 = ~pi26 & n4071;
  assign n4073 = ~n3785 & ~n4026;
  assign n4074 = n3785 & n4026;
  assign n4075 = ~n4073 & ~n4074;
  assign n4076 = ~n3973 & ~n4075;
  assign n4077 = ~n3782 & n3973;
  assign n4078 = ~n4076 & ~n4077;
  assign n4079 = pi21 & n4078;
  assign n4080 = ~pi21 & ~n4078;
  assign n4081 = ~n4079 & ~n4080;
  assign n4082 = ~n3730 & ~n4024;
  assign n4083 = n3730 & n4024;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~n3973 & ~n4084;
  assign n4086 = n3727 & n3973;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = ~pi20 & ~n4087;
  assign n4089 = pi20 & n4087;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = n4072 & n4090;
  assign n4092 = n4081 & n4091;
  assign n4093 = n4069 & n4092;
  assign n4094 = n4049 & n4093;
  assign n4095 = n4040 & n4094;
  assign n4096 = n4060 & n4095;
  assign n4097 = ~n3800 & ~n4022;
  assign n4098 = n3800 & n4022;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = ~n3973 & ~n4099;
  assign n4101 = ~n3797 & n3973;
  assign n4102 = ~n4100 & ~n4101;
  assign n4103 = pi19 & n4102;
  assign n4104 = ~pi19 & ~n4102;
  assign n4105 = ~n4103 & ~n4104;
  assign n4106 = n3815 & n3973;
  assign n4107 = ~n3818 & ~n4018;
  assign n4108 = n3818 & n4018;
  assign n4109 = ~n3973 & ~n4107;
  assign n4110 = ~n4108 & n4109;
  assign n4111 = ~n4106 & ~n4110;
  assign n4112 = pi17 & n4111;
  assign n4113 = ~pi17 & ~n4111;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = ~n3806 & n3973;
  assign n4116 = n3809 & ~n4016;
  assign n4117 = ~n3809 & n4016;
  assign n4118 = ~n3973 & ~n4116;
  assign n4119 = ~n4117 & n4118;
  assign n4120 = ~n4115 & ~n4119;
  assign n4121 = pi16 & ~n4120;
  assign n4122 = ~pi16 & n4120;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = ~n3824 & n3973;
  assign n4125 = n3827 & ~n4020;
  assign n4126 = ~n3827 & n4020;
  assign n4127 = ~n3973 & ~n4125;
  assign n4128 = ~n4126 & n4127;
  assign n4129 = ~n4124 & ~n4128;
  assign n4130 = pi18 & ~n4129;
  assign n4131 = ~pi18 & n4129;
  assign n4132 = ~n4130 & ~n4131;
  assign n4133 = n4114 & n4123;
  assign n4134 = n4132 & n4133;
  assign n4135 = n4105 & n4134;
  assign n4136 = n4096 & n4135;
  assign n4137 = ~n3866 & n3973;
  assign n4138 = n3869 & ~n4014;
  assign n4139 = ~n3869 & n4014;
  assign n4140 = ~n4138 & ~n4139;
  assign n4141 = ~n3973 & n4140;
  assign n4142 = ~n4137 & ~n4141;
  assign n4143 = pi15 & ~n4142;
  assign n4144 = ~pi15 & n4142;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = ~n3847 & n3973;
  assign n4147 = n3850 & ~n4008;
  assign n4148 = ~n3850 & n4008;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = ~n3973 & n4149;
  assign n4151 = ~n4146 & ~n4150;
  assign n4152 = pi12 & n4151;
  assign n4153 = ~pi12 & ~n4151;
  assign n4154 = ~n4152 & ~n4153;
  assign n4155 = n3838 & n3973;
  assign n4156 = n3841 & ~n4010;
  assign n4157 = ~n3841 & n4010;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = ~n3973 & n4158;
  assign n4160 = ~n4155 & ~n4159;
  assign n4161 = pi13 & n4160;
  assign n4162 = ~pi13 & ~n4160;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = ~n3857 & n3973;
  assign n4165 = n3860 & ~n4012;
  assign n4166 = ~n3860 & n4012;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = ~n3973 & n4167;
  assign n4169 = ~n4164 & ~n4168;
  assign n4170 = pi14 & ~n4169;
  assign n4171 = ~pi14 & n4169;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = n4145 & n4154;
  assign n4174 = n4163 & n4172;
  assign n4175 = n4173 & n4174;
  assign n4176 = n4136 & n4175;
  assign n4177 = ~n3674 & n3973;
  assign n4178 = n3940 & ~n4006;
  assign n4179 = ~n3940 & n4006;
  assign n4180 = ~n4178 & ~n4179;
  assign n4181 = ~n3973 & n4180;
  assign n4182 = ~n4177 & ~n4181;
  assign n4183 = ~pi11 & ~n4182;
  assign n4184 = pi11 & n4182;
  assign n4185 = ~n4183 & ~n4184;
  assign n4186 = ~n3941 & ~n4004;
  assign n4187 = n3941 & n4004;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~n3973 & ~n4188;
  assign n4190 = ~n3682 & n3973;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = ~pi10 & ~n4191;
  assign n4193 = pi10 & n4191;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = n3689 & n3973;
  assign n4196 = n3942 & ~n4002;
  assign n4197 = ~n3942 & n4002;
  assign n4198 = ~n4196 & ~n4197;
  assign n4199 = ~n3973 & n4198;
  assign n4200 = ~n4195 & ~n4199;
  assign n4201 = pi09 & ~n4200;
  assign n4202 = ~pi09 & n4200;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = ~n3696 & n3973;
  assign n4205 = n3944 & ~n4000;
  assign n4206 = ~n3944 & n4000;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = ~n3973 & n4207;
  assign n4209 = ~n4204 & ~n4208;
  assign n4210 = pi08 & ~n4209;
  assign n4211 = ~pi08 & n4209;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = n4185 & n4194;
  assign n4214 = n4203 & n4212;
  assign n4215 = n4213 & n4214;
  assign n4216 = n4176 & n4215;
  assign n4217 = ~n3931 & n3973;
  assign n4218 = n3955 & ~n3983;
  assign n4219 = ~n3955 & n3983;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = ~n3973 & n4220;
  assign n4222 = ~n4217 & ~n4221;
  assign n4223 = ~pi04 & ~n4222;
  assign n4224 = pi04 & n4222;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = n3924 & n3973;
  assign n4227 = n3953 & ~n3985;
  assign n4228 = ~n3953 & n3985;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n3973 & n4229;
  assign n4231 = ~n4226 & ~n4230;
  assign n4232 = ~pi05 & ~n4231;
  assign n4233 = pi05 & n4231;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = ~n3909 & n3973;
  assign n4236 = ~n3952 & ~n3998;
  assign n4237 = n3952 & n3998;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = ~n3973 & n4238;
  assign n4240 = ~n4235 & ~n4239;
  assign n4241 = pi07 & ~n4240;
  assign n4242 = ~pi07 & n4240;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = n3995 & n4225;
  assign n4245 = n4234 & n4243;
  assign n4246 = n4244 & n4245;
  assign n4247 = n4216 & n4246;
  assign n4248 = ~pi03 & n3980;
  assign n4249 = pi03 & ~n3980;
  assign n4250 = pi00 & ~n3639;
  assign n4251 = n3642 & n3652;
  assign n4252 = ~pi01 & ~n4251;
  assign n4253 = n4250 & n4252;
  assign n4254 = pi01 & ~n4250;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = ~n3973 & n4255;
  assign n4257 = ~n3964 & n3973;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = pi02 & ~n4258;
  assign n4260 = ~n4249 & ~n4259;
  assign n4261 = ~n4248 & ~n4260;
  assign n4262 = n4247 & ~n4261;
  assign n4263 = n4153 & ~n4161;
  assign n4264 = ~n4162 & ~n4171;
  assign n4265 = ~n4263 & n4264;
  assign n4266 = ~n4143 & ~n4170;
  assign n4267 = ~n4265 & n4266;
  assign n4268 = ~n4144 & ~n4267;
  assign n4269 = n4136 & n4268;
  assign n4270 = ~n4113 & n4121;
  assign n4271 = ~n4112 & ~n4270;
  assign n4272 = ~n4130 & n4271;
  assign n4273 = ~n4131 & ~n4272;
  assign n4274 = ~n4104 & n4273;
  assign n4275 = ~n4103 & ~n4274;
  assign n4276 = n4096 & n4275;
  assign n4277 = ~n4080 & ~n4088;
  assign n4278 = ~n4079 & ~n4277;
  assign n4279 = ~n4067 & n4278;
  assign n4280 = ~n4068 & ~n4279;
  assign n4281 = ~n4048 & n4280;
  assign n4282 = ~n4047 & ~n4281;
  assign n4283 = ~n4038 & n4282;
  assign n4284 = ~n4039 & ~n4283;
  assign n4285 = ~n4059 & n4284;
  assign n4286 = ~n4058 & n4072;
  assign n4287 = ~n4285 & n4286;
  assign n4288 = ~n4276 & ~n4287;
  assign n4289 = ~n4269 & ~n4288;
  assign n4290 = ~n4202 & n4210;
  assign n4291 = ~n4193 & ~n4201;
  assign n4292 = ~n4290 & n4291;
  assign n4293 = ~n4183 & ~n4192;
  assign n4294 = ~n4292 & n4293;
  assign n4295 = ~n4184 & ~n4294;
  assign n4296 = n4176 & n4295;
  assign n4297 = ~n4216 & ~n4289;
  assign n4298 = ~n4296 & n4297;
  assign n4299 = ~n4223 & ~n4232;
  assign n4300 = ~n3993 & ~n4233;
  assign n4301 = ~n4299 & n4300;
  assign n4302 = ~n3994 & ~n4301;
  assign n4303 = ~n4241 & ~n4302;
  assign n4304 = ~n4242 & ~n4303;
  assign n4305 = n4216 & n4304;
  assign n4306 = ~n4298 & ~n4305;
  assign n4307 = ~n4262 & ~n4306;
  assign n4308 = ~pi02 & n4258;
  assign n4309 = ~n4259 & ~n4308;
  assign n4310 = ~n4248 & ~n4249;
  assign n4311 = n4309 & n4310;
  assign n4312 = n4247 & n4311;
  assign n4313 = ~n4307 & ~n4312;
  assign n4314 = pi00 & n3973;
  assign n4315 = ~pi01 & ~n4314;
  assign n4316 = n4312 & n4315;
  assign n4317 = ~n4313 & ~n4316;
  assign n4318 = ~n3980 & n4317;
  assign n4319 = ~n4308 & ~n4315;
  assign n4320 = ~n4259 & ~n4319;
  assign n4321 = n4310 & ~n4320;
  assign n4322 = ~n4310 & n4320;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = ~n4317 & n4323;
  assign n4325 = ~n4318 & ~n4324;
  assign n4326 = pi04 & ~n4325;
  assign n4327 = ~pi04 & n4325;
  assign n4328 = n4258 & n4317;
  assign n4329 = ~n4309 & ~n4315;
  assign n4330 = n4309 & n4315;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = ~n4317 & n4331;
  assign n4333 = ~n4328 & ~n4332;
  assign n4334 = pi03 & n4333;
  assign n4335 = pi00 & ~n3969;
  assign n4336 = ~pi01 & ~n4335;
  assign n4337 = pi01 & n4335;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = ~n4317 & ~n4338;
  assign n4340 = pi00 & ~n3973;
  assign n4341 = n4317 & ~n4340;
  assign n4342 = ~n4339 & ~n4341;
  assign n4343 = ~pi02 & n4342;
  assign n4344 = pi02 & ~n4342;
  assign n4345 = pi00 & ~n4317;
  assign n4346 = ~pi01 & n4345;
  assign n4347 = ~n4344 & n4346;
  assign n4348 = ~pi03 & ~n4333;
  assign n4349 = ~n4343 & ~n4348;
  assign n4350 = ~n4347 & n4349;
  assign n4351 = ~n4334 & ~n4350;
  assign n4352 = ~n4327 & ~n4351;
  assign n4353 = ~n4249 & n4320;
  assign n4354 = ~n4248 & ~n4353;
  assign n4355 = ~n4224 & ~n4354;
  assign n4356 = ~n4223 & ~n4355;
  assign n4357 = ~n4232 & n4356;
  assign n4358 = ~n4233 & ~n4357;
  assign n4359 = ~n3993 & n4358;
  assign n4360 = ~n3994 & ~n4359;
  assign n4361 = ~n4242 & n4360;
  assign n4362 = ~n4241 & ~n4361;
  assign n4363 = ~n4211 & ~n4362;
  assign n4364 = ~n4210 & ~n4363;
  assign n4365 = ~n4202 & ~n4364;
  assign n4366 = ~n4201 & ~n4365;
  assign n4367 = ~n4192 & ~n4366;
  assign n4368 = ~n4193 & ~n4367;
  assign n4369 = ~n4183 & ~n4368;
  assign n4370 = ~n4184 & ~n4369;
  assign n4371 = ~n4152 & n4370;
  assign n4372 = ~n4153 & ~n4371;
  assign n4373 = ~n4161 & ~n4372;
  assign n4374 = ~n4162 & ~n4373;
  assign n4375 = ~n4171 & n4374;
  assign n4376 = ~n4170 & ~n4375;
  assign n4377 = ~n4144 & ~n4376;
  assign n4378 = ~n4143 & ~n4377;
  assign n4379 = ~n4122 & ~n4378;
  assign n4380 = ~n4121 & ~n4379;
  assign n4381 = ~n4112 & n4380;
  assign n4382 = ~n4113 & ~n4381;
  assign n4383 = ~n4130 & ~n4382;
  assign n4384 = ~n4131 & ~n4383;
  assign n4385 = ~n4103 & ~n4384;
  assign n4386 = ~n4104 & ~n4385;
  assign n4387 = ~n4089 & ~n4386;
  assign n4388 = ~n4088 & ~n4387;
  assign n4389 = ~n4079 & ~n4388;
  assign n4390 = ~n4080 & ~n4389;
  assign n4391 = ~n4067 & ~n4390;
  assign n4392 = ~n4068 & ~n4391;
  assign n4393 = ~n4049 & ~n4392;
  assign n4394 = n4049 & n4392;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = ~n4317 & ~n4395;
  assign n4397 = ~n4046 & n4317;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = pi24 & n4398;
  assign n4400 = ~pi24 & ~n4398;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = ~n4090 & ~n4386;
  assign n4403 = n4090 & n4386;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4317 & ~n4404;
  assign n4406 = ~n4087 & n4317;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = ~pi21 & ~n4407;
  assign n4409 = ~n4081 & ~n4388;
  assign n4410 = n4081 & n4388;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4317 & ~n4411;
  assign n4413 = ~n4078 & n4317;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = pi22 & n4414;
  assign n4416 = ~pi22 & ~n4414;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418 = ~n4066 & n4317;
  assign n4419 = n4069 & ~n4390;
  assign n4420 = ~n4069 & n4390;
  assign n4421 = ~n4317 & ~n4419;
  assign n4422 = ~n4420 & n4421;
  assign n4423 = ~n4418 & ~n4422;
  assign n4424 = pi23 & n4423;
  assign n4425 = ~pi23 & ~n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = n4071 & ~n4408;
  assign n4428 = n4417 & n4427;
  assign n4429 = n4426 & n4428;
  assign n4430 = ~n4057 & n4317;
  assign n4431 = ~n4047 & ~n4392;
  assign n4432 = ~n4048 & ~n4431;
  assign n4433 = ~n4039 & n4432;
  assign n4434 = ~n4038 & ~n4433;
  assign n4435 = n4060 & ~n4434;
  assign n4436 = ~n4060 & n4434;
  assign n4437 = ~n4317 & ~n4435;
  assign n4438 = ~n4436 & n4437;
  assign n4439 = ~n4430 & ~n4438;
  assign n4440 = pi26 & ~n4439;
  assign n4441 = ~pi26 & n4439;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~n4037 & n4317;
  assign n4444 = ~n4040 & ~n4432;
  assign n4445 = n4040 & n4432;
  assign n4446 = ~n4317 & ~n4444;
  assign n4447 = ~n4445 & n4446;
  assign n4448 = ~n4443 & ~n4447;
  assign n4449 = pi25 & ~n4448;
  assign n4450 = ~pi25 & n4448;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = pi21 & n4407;
  assign n4453 = n4429 & ~n4452;
  assign n4454 = n4401 & n4453;
  assign n4455 = n4451 & n4454;
  assign n4456 = n4442 & n4455;
  assign n4457 = ~n4105 & ~n4384;
  assign n4458 = n4105 & n4384;
  assign n4459 = ~n4457 & ~n4458;
  assign n4460 = ~n4317 & ~n4459;
  assign n4461 = ~n4102 & n4317;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = pi20 & n4462;
  assign n4464 = ~pi20 & ~n4462;
  assign n4465 = ~n4463 & ~n4464;
  assign n4466 = ~n4123 & ~n4378;
  assign n4467 = n4123 & n4378;
  assign n4468 = ~n4466 & ~n4467;
  assign n4469 = ~n4317 & ~n4468;
  assign n4470 = ~n4120 & n4317;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = pi17 & ~n4471;
  assign n4473 = ~pi17 & n4471;
  assign n4474 = ~n4472 & ~n4473;
  assign n4475 = n4111 & n4317;
  assign n4476 = n4114 & ~n4380;
  assign n4477 = ~n4114 & n4380;
  assign n4478 = ~n4317 & ~n4476;
  assign n4479 = ~n4477 & n4478;
  assign n4480 = ~n4475 & ~n4479;
  assign n4481 = pi18 & ~n4480;
  assign n4482 = ~pi18 & n4480;
  assign n4483 = ~n4481 & ~n4482;
  assign n4484 = n4129 & n4317;
  assign n4485 = n4132 & ~n4382;
  assign n4486 = ~n4132 & n4382;
  assign n4487 = ~n4317 & ~n4485;
  assign n4488 = ~n4486 & n4487;
  assign n4489 = ~n4484 & ~n4488;
  assign n4490 = pi19 & n4489;
  assign n4491 = ~pi19 & ~n4489;
  assign n4492 = ~n4490 & ~n4491;
  assign n4493 = n4474 & n4483;
  assign n4494 = n4492 & n4493;
  assign n4495 = n4465 & n4494;
  assign n4496 = n4456 & n4495;
  assign n4497 = ~n4160 & n4317;
  assign n4498 = n4163 & ~n4372;
  assign n4499 = ~n4163 & n4372;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = ~n4317 & n4500;
  assign n4502 = ~n4497 & ~n4501;
  assign n4503 = pi14 & n4502;
  assign n4504 = ~pi14 & ~n4502;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = ~n4145 & ~n4376;
  assign n4507 = n4145 & n4376;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = ~n4317 & ~n4508;
  assign n4510 = ~n4142 & n4317;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = pi16 & ~n4511;
  assign n4513 = ~pi16 & n4511;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = n4151 & n4317;
  assign n4516 = n4154 & ~n4370;
  assign n4517 = ~n4154 & n4370;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = ~n4317 & n4518;
  assign n4520 = ~n4515 & ~n4519;
  assign n4521 = pi13 & ~n4520;
  assign n4522 = ~pi13 & n4520;
  assign n4523 = ~n4521 & ~n4522;
  assign n4524 = n4169 & n4317;
  assign n4525 = n4172 & ~n4374;
  assign n4526 = ~n4172 & n4374;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = ~n4317 & n4527;
  assign n4529 = ~n4524 & ~n4528;
  assign n4530 = pi15 & n4529;
  assign n4531 = ~pi15 & ~n4529;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = n4505 & n4514;
  assign n4534 = n4523 & n4532;
  assign n4535 = n4533 & n4534;
  assign n4536 = n4496 & n4535;
  assign n4537 = n4182 & n4317;
  assign n4538 = n4185 & ~n4368;
  assign n4539 = ~n4185 & n4368;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = ~n4317 & n4540;
  assign n4542 = ~n4537 & ~n4541;
  assign n4543 = pi12 & ~n4542;
  assign n4544 = ~pi12 & n4542;
  assign n4545 = ~n4543 & ~n4544;
  assign n4546 = n4191 & n4317;
  assign n4547 = n4194 & ~n4366;
  assign n4548 = ~n4194 & n4366;
  assign n4549 = ~n4547 & ~n4548;
  assign n4550 = ~n4317 & n4549;
  assign n4551 = ~n4546 & ~n4550;
  assign n4552 = pi11 & ~n4551;
  assign n4553 = ~pi11 & n4551;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = ~n4200 & n4317;
  assign n4556 = n4203 & ~n4364;
  assign n4557 = ~n4203 & n4364;
  assign n4558 = ~n4556 & ~n4557;
  assign n4559 = ~n4317 & n4558;
  assign n4560 = ~n4555 & ~n4559;
  assign n4561 = pi10 & ~n4560;
  assign n4562 = ~pi10 & n4560;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = ~n4209 & n4317;
  assign n4565 = n4212 & ~n4362;
  assign n4566 = ~n4212 & n4362;
  assign n4567 = ~n4565 & ~n4566;
  assign n4568 = ~n4317 & n4567;
  assign n4569 = ~n4564 & ~n4568;
  assign n4570 = pi09 & ~n4569;
  assign n4571 = ~pi09 & n4569;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4545 & n4554;
  assign n4574 = n4563 & n4572;
  assign n4575 = n4573 & n4574;
  assign n4576 = n4536 & n4575;
  assign n4577 = n3992 & n4317;
  assign n4578 = ~n3995 & ~n4358;
  assign n4579 = n3995 & n4358;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~n4317 & n4580;
  assign n4582 = ~n4577 & ~n4581;
  assign n4583 = pi07 & n4582;
  assign n4584 = ~pi07 & ~n4582;
  assign n4585 = ~n4583 & ~n4584;
  assign n4586 = ~n4231 & n4317;
  assign n4587 = n4234 & ~n4356;
  assign n4588 = ~n4234 & n4356;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = ~n4317 & n4589;
  assign n4591 = ~n4586 & ~n4590;
  assign n4592 = pi06 & n4591;
  assign n4593 = ~pi06 & ~n4591;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = ~n4225 & ~n4354;
  assign n4596 = n4225 & n4354;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = ~n4317 & ~n4597;
  assign n4599 = ~n4222 & n4317;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = pi05 & n4600;
  assign n4602 = ~pi05 & ~n4600;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = ~n4240 & n4317;
  assign n4605 = ~n4243 & ~n4360;
  assign n4606 = n4243 & n4360;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4317 & n4607;
  assign n4609 = ~n4604 & ~n4608;
  assign n4610 = pi08 & ~n4609;
  assign n4611 = ~pi08 & n4609;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = n4585 & n4594;
  assign n4614 = n4603 & n4612;
  assign n4615 = n4613 & n4614;
  assign n4616 = n4576 & n4615;
  assign n4617 = ~n4326 & ~n4352;
  assign n4618 = n4616 & n4617;
  assign n4619 = n4472 & ~n4482;
  assign n4620 = ~n4481 & ~n4619;
  assign n4621 = ~n4490 & n4620;
  assign n4622 = ~n4491 & ~n4621;
  assign n4623 = ~n4464 & n4622;
  assign n4624 = ~n4463 & ~n4623;
  assign n4625 = n4456 & n4624;
  assign n4626 = ~n4415 & ~n4424;
  assign n4627 = ~n4425 & ~n4626;
  assign n4628 = ~n4399 & ~n4429;
  assign n4629 = ~n4627 & n4628;
  assign n4630 = ~n4400 & ~n4450;
  assign n4631 = ~n4629 & n4630;
  assign n4632 = ~n4440 & ~n4449;
  assign n4633 = ~n4631 & n4632;
  assign n4634 = ~n4441 & ~n4633;
  assign n4635 = n4071 & ~n4634;
  assign n4636 = ~n4625 & ~n4635;
  assign n4637 = ~n4503 & n4522;
  assign n4638 = ~n4504 & ~n4531;
  assign n4639 = ~n4637 & n4638;
  assign n4640 = ~n4512 & ~n4530;
  assign n4641 = ~n4639 & n4640;
  assign n4642 = ~n4513 & ~n4641;
  assign n4643 = n4496 & n4642;
  assign n4644 = ~n4636 & ~n4643;
  assign n4645 = ~n4561 & ~n4570;
  assign n4646 = ~n4553 & ~n4562;
  assign n4647 = ~n4645 & n4646;
  assign n4648 = ~n4543 & ~n4552;
  assign n4649 = ~n4647 & n4648;
  assign n4650 = ~n4544 & ~n4649;
  assign n4651 = n4536 & ~n4650;
  assign n4652 = ~n4644 & ~n4651;
  assign n4653 = ~n4593 & ~n4602;
  assign n4654 = ~n4583 & ~n4592;
  assign n4655 = ~n4653 & n4654;
  assign n4656 = ~n4584 & ~n4611;
  assign n4657 = ~n4655 & n4656;
  assign n4658 = ~n4610 & ~n4657;
  assign n4659 = n4576 & ~n4658;
  assign n4660 = ~n4652 & ~n4659;
  assign n4661 = ~n4618 & ~n4660;
  assign n4662 = ~n4343 & ~n4344;
  assign n4663 = ~n4326 & ~n4327;
  assign n4664 = ~n4334 & ~n4348;
  assign n4665 = n84 & n4662;
  assign n4666 = n4663 & n4664;
  assign n4667 = n4665 & n4666;
  assign n4668 = n4616 & n4667;
  assign n4669 = n4661 & ~n4668;
  assign n4670 = ~n84 & ~n4346;
  assign n4671 = ~n4343 & n4670;
  assign n4672 = ~n4344 & ~n4671;
  assign n4673 = ~n4348 & ~n4672;
  assign n4674 = ~n4334 & ~n4673;
  assign n4675 = ~n4327 & ~n4674;
  assign n4676 = ~n4326 & ~n4675;
  assign n4677 = ~n4601 & n4676;
  assign n4678 = ~n4602 & ~n4677;
  assign n4679 = ~n4593 & n4678;
  assign n4680 = ~n4592 & ~n4679;
  assign n4681 = ~n4584 & ~n4680;
  assign n4682 = ~n4583 & ~n4681;
  assign n4683 = ~n4610 & n4682;
  assign n4684 = ~n4611 & ~n4683;
  assign n4685 = ~n4570 & ~n4684;
  assign n4686 = ~n4571 & ~n4685;
  assign n4687 = ~n4562 & n4686;
  assign n4688 = ~n4561 & ~n4687;
  assign n4689 = ~n4553 & ~n4688;
  assign n4690 = ~n4552 & ~n4689;
  assign n4691 = ~n4543 & n4690;
  assign n4692 = ~n4544 & ~n4691;
  assign n4693 = ~n4523 & ~n4692;
  assign n4694 = n4523 & n4692;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4669 & ~n4695;
  assign n4697 = n4520 & n4669;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = n4600 & n4669;
  assign n4700 = n4603 & ~n4676;
  assign n4701 = ~n4603 & n4676;
  assign n4702 = ~n4700 & ~n4701;
  assign n4703 = ~n4669 & n4702;
  assign n4704 = ~n4699 & ~n4703;
  assign n4705 = pi06 & ~n4704;
  assign n4706 = ~n4594 & ~n4678;
  assign n4707 = n4594 & n4678;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n4669 & ~n4708;
  assign n4710 = ~n4591 & n4669;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = pi07 & n4711;
  assign n4713 = ~pi07 & ~n4711;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = ~n4609 & n4669;
  assign n4716 = n4612 & ~n4682;
  assign n4717 = ~n4612 & n4682;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = ~n4669 & n4718;
  assign n4720 = ~n4715 & ~n4719;
  assign n4721 = pi09 & ~n4720;
  assign n4722 = ~pi09 & n4720;
  assign n4723 = ~n4721 & ~n4722;
  assign n4724 = ~pi06 & n4704;
  assign n4725 = ~n4585 & ~n4680;
  assign n4726 = n4585 & n4680;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = ~n4669 & ~n4727;
  assign n4729 = n4582 & n4669;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = pi08 & ~n4730;
  assign n4732 = ~pi08 & n4730;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = n4714 & ~n4724;
  assign n4735 = n4723 & n4733;
  assign n4736 = n4734 & n4735;
  assign n4737 = pi14 & n4698;
  assign n4738 = n4407 & n4669;
  assign n4739 = ~n4408 & ~n4452;
  assign n4740 = ~n4521 & ~n4692;
  assign n4741 = ~n4522 & ~n4740;
  assign n4742 = ~n4503 & ~n4741;
  assign n4743 = ~n4504 & ~n4742;
  assign n4744 = ~n4530 & ~n4743;
  assign n4745 = ~n4531 & ~n4744;
  assign n4746 = ~n4512 & ~n4745;
  assign n4747 = ~n4513 & ~n4746;
  assign n4748 = ~n4473 & n4747;
  assign n4749 = ~n4472 & ~n4748;
  assign n4750 = ~n4482 & ~n4749;
  assign n4751 = ~n4481 & ~n4750;
  assign n4752 = ~n4490 & n4751;
  assign n4753 = ~n4491 & ~n4752;
  assign n4754 = ~n4463 & ~n4753;
  assign n4755 = ~n4464 & ~n4754;
  assign n4756 = ~n4739 & ~n4755;
  assign n4757 = n4739 & n4755;
  assign n4758 = ~n4669 & ~n4756;
  assign n4759 = ~n4757 & n4758;
  assign n4760 = ~n4738 & ~n4759;
  assign n4761 = pi22 & ~n4760;
  assign n4762 = ~n4452 & ~n4755;
  assign n4763 = ~n4408 & ~n4762;
  assign n4764 = ~n4415 & ~n4763;
  assign n4765 = ~n4416 & ~n4764;
  assign n4766 = ~n4426 & ~n4765;
  assign n4767 = n4426 & n4765;
  assign n4768 = ~n4766 & ~n4767;
  assign n4769 = ~n4669 & ~n4768;
  assign n4770 = ~n4423 & n4669;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = pi24 & n4771;
  assign n4773 = ~pi24 & ~n4771;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = ~n4398 & n4669;
  assign n4776 = ~n4424 & ~n4765;
  assign n4777 = ~n4425 & ~n4776;
  assign n4778 = n4401 & ~n4777;
  assign n4779 = ~n4401 & n4777;
  assign n4780 = ~n4669 & ~n4778;
  assign n4781 = ~n4779 & n4780;
  assign n4782 = ~n4775 & ~n4781;
  assign n4783 = pi25 & n4782;
  assign n4784 = ~pi25 & ~n4782;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~n4439 & n4669;
  assign n4787 = ~n4399 & ~n4777;
  assign n4788 = ~n4400 & ~n4787;
  assign n4789 = ~n4449 & ~n4788;
  assign n4790 = ~n4450 & ~n4789;
  assign n4791 = ~n4442 & ~n4790;
  assign n4792 = n4442 & n4790;
  assign n4793 = ~n4669 & ~n4791;
  assign n4794 = ~n4792 & n4793;
  assign n4795 = ~n4786 & ~n4794;
  assign n4796 = pi27 & ~n4795;
  assign n4797 = ~pi27 & n4795;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~n4451 & ~n4788;
  assign n4800 = n4451 & n4788;
  assign n4801 = ~n4799 & ~n4800;
  assign n4802 = ~n4669 & ~n4801;
  assign n4803 = n4448 & n4669;
  assign n4804 = ~n4802 & ~n4803;
  assign n4805 = pi26 & n4804;
  assign n4806 = ~pi26 & ~n4804;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = ~pi22 & n4760;
  assign n4809 = ~n4417 & ~n4763;
  assign n4810 = n4417 & n4763;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = ~n4669 & ~n4811;
  assign n4813 = ~n4414 & n4669;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = pi23 & n4814;
  assign n4816 = ~pi23 & ~n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n4070 & ~n4808;
  assign n4819 = n4817 & n4818;
  assign n4820 = n4774 & n4819;
  assign n4821 = n4785 & n4820;
  assign n4822 = n4807 & n4821;
  assign n4823 = n4798 & n4822;
  assign n4824 = ~n4761 & n4823;
  assign n4825 = ~n4465 & ~n4753;
  assign n4826 = n4465 & n4753;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n4669 & ~n4827;
  assign n4829 = ~n4462 & n4669;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = pi21 & n4830;
  assign n4832 = ~pi21 & ~n4830;
  assign n4833 = ~n4831 & ~n4832;
  assign n4834 = n4471 & n4669;
  assign n4835 = n4474 & ~n4747;
  assign n4836 = ~n4474 & n4747;
  assign n4837 = ~n4669 & ~n4835;
  assign n4838 = ~n4836 & n4837;
  assign n4839 = ~n4834 & ~n4838;
  assign n4840 = pi18 & n4839;
  assign n4841 = ~pi18 & ~n4839;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~n4480 & n4669;
  assign n4844 = n4483 & ~n4749;
  assign n4845 = ~n4483 & n4749;
  assign n4846 = ~n4669 & ~n4844;
  assign n4847 = ~n4845 & n4846;
  assign n4848 = ~n4843 & ~n4847;
  assign n4849 = pi19 & ~n4848;
  assign n4850 = ~pi19 & n4848;
  assign n4851 = ~n4849 & ~n4850;
  assign n4852 = ~n4492 & ~n4751;
  assign n4853 = n4492 & n4751;
  assign n4854 = ~n4852 & ~n4853;
  assign n4855 = ~n4669 & ~n4854;
  assign n4856 = n4489 & n4669;
  assign n4857 = ~n4855 & ~n4856;
  assign n4858 = pi20 & ~n4857;
  assign n4859 = ~pi20 & n4857;
  assign n4860 = ~n4858 & ~n4859;
  assign n4861 = n4842 & n4851;
  assign n4862 = n4860 & n4861;
  assign n4863 = n4833 & n4862;
  assign n4864 = n4824 & n4863;
  assign n4865 = ~n4514 & ~n4745;
  assign n4866 = n4514 & n4745;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n4669 & ~n4867;
  assign n4869 = n4511 & n4669;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = pi17 & n4870;
  assign n4872 = ~pi17 & ~n4870;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = ~n4529 & n4669;
  assign n4875 = n4532 & ~n4743;
  assign n4876 = ~n4532 & n4743;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = ~n4669 & n4877;
  assign n4879 = ~n4874 & ~n4878;
  assign n4880 = pi16 & n4879;
  assign n4881 = ~pi16 & ~n4879;
  assign n4882 = ~n4880 & ~n4881;
  assign n4883 = ~pi14 & ~n4698;
  assign n4884 = ~n4505 & ~n4741;
  assign n4885 = n4505 & n4741;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = ~n4669 & ~n4886;
  assign n4888 = ~n4502 & n4669;
  assign n4889 = ~n4887 & ~n4888;
  assign n4890 = pi15 & n4889;
  assign n4891 = ~pi15 & ~n4889;
  assign n4892 = ~n4890 & ~n4891;
  assign n4893 = n4882 & ~n4883;
  assign n4894 = n4892 & n4893;
  assign n4895 = n4873 & n4894;
  assign n4896 = ~n4737 & n4895;
  assign n4897 = n4864 & n4896;
  assign n4898 = ~n4542 & n4669;
  assign n4899 = n4545 & ~n4690;
  assign n4900 = ~n4545 & n4690;
  assign n4901 = ~n4899 & ~n4900;
  assign n4902 = ~n4669 & n4901;
  assign n4903 = ~n4898 & ~n4902;
  assign n4904 = pi13 & ~n4903;
  assign n4905 = ~pi13 & n4903;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = ~n4551 & n4669;
  assign n4908 = n4554 & ~n4688;
  assign n4909 = ~n4554 & n4688;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = ~n4669 & n4910;
  assign n4912 = ~n4907 & ~n4911;
  assign n4913 = pi12 & ~n4912;
  assign n4914 = ~pi12 & n4912;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = ~n4560 & n4669;
  assign n4917 = ~n4563 & ~n4686;
  assign n4918 = n4563 & n4686;
  assign n4919 = ~n4917 & ~n4918;
  assign n4920 = ~n4669 & n4919;
  assign n4921 = ~n4916 & ~n4920;
  assign n4922 = pi11 & ~n4921;
  assign n4923 = ~pi11 & n4921;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = ~n4572 & ~n4684;
  assign n4926 = n4572 & n4684;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 = ~n4669 & ~n4927;
  assign n4929 = n4569 & n4669;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = pi10 & n4930;
  assign n4932 = ~pi10 & ~n4930;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = n4906 & n4915;
  assign n4935 = n4924 & n4933;
  assign n4936 = n4934 & n4935;
  assign n4937 = n4897 & n4936;
  assign n4938 = ~n4705 & n4736;
  assign n4939 = n4937 & n4938;
  assign n4940 = ~n4325 & n4669;
  assign n4941 = n4663 & ~n4674;
  assign n4942 = ~n4663 & n4674;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4669 & n4943;
  assign n4945 = ~n4940 & ~n4944;
  assign n4946 = pi05 & ~n4945;
  assign n4947 = n4333 & n4669;
  assign n4948 = n4664 & ~n4672;
  assign n4949 = ~n4664 & n4672;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4669 & n4950;
  assign n4952 = ~n4947 & ~n4951;
  assign n4953 = ~pi04 & n4952;
  assign n4954 = ~pi05 & n4945;
  assign n4955 = ~n4342 & n4669;
  assign n4956 = ~n4662 & ~n4670;
  assign n4957 = n4662 & n4670;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4669 & n4958;
  assign n4960 = ~n4955 & ~n4959;
  assign n4961 = pi03 & ~n4960;
  assign n4962 = pi04 & ~n4952;
  assign n4963 = ~pi03 & n4960;
  assign n4964 = pi00 & ~n4313;
  assign n4965 = n4312 & n4340;
  assign n4966 = ~pi01 & ~n4965;
  assign n4967 = n4964 & n4966;
  assign n4968 = pi01 & ~n4964;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = ~n4669 & n4969;
  assign n4971 = ~n4345 & n4669;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = pi02 & ~n4972;
  assign n4974 = ~n4963 & n4973;
  assign n4975 = ~n4961 & ~n4962;
  assign n4976 = ~n4974 & n4975;
  assign n4977 = ~n4953 & ~n4954;
  assign n4978 = ~n4976 & n4977;
  assign n4979 = ~n4946 & ~n4978;
  assign n4980 = n4939 & n4979;
  assign n4981 = ~n4773 & n4815;
  assign n4982 = ~n4772 & ~n4981;
  assign n4983 = ~n4783 & n4982;
  assign n4984 = ~n4784 & ~n4983;
  assign n4985 = ~n4806 & n4984;
  assign n4986 = ~n4805 & ~n4985;
  assign n4987 = ~n4797 & ~n4986;
  assign n4988 = n4070 & ~n4796;
  assign n4989 = ~n4987 & n4988;
  assign n4990 = ~n4823 & n4989;
  assign n4991 = n4840 & ~n4850;
  assign n4992 = ~n4849 & ~n4991;
  assign n4993 = ~n4858 & n4992;
  assign n4994 = ~n4859 & ~n4993;
  assign n4995 = ~n4832 & n4994;
  assign n4996 = ~n4831 & ~n4995;
  assign n4997 = n4824 & n4996;
  assign n4998 = ~n4864 & ~n4990;
  assign n4999 = ~n4997 & n4998;
  assign n5000 = ~n4880 & ~n4890;
  assign n5001 = ~n4881 & ~n5000;
  assign n5002 = ~n4872 & n5001;
  assign n5003 = ~n4871 & ~n5002;
  assign n5004 = ~n4895 & n5003;
  assign n5005 = n4864 & ~n5004;
  assign n5006 = ~n4999 & ~n5005;
  assign n5007 = ~n4922 & ~n4931;
  assign n5008 = ~n4914 & ~n4923;
  assign n5009 = ~n5007 & n5008;
  assign n5010 = ~n4904 & ~n4913;
  assign n5011 = ~n5009 & n5010;
  assign n5012 = ~n4905 & ~n5011;
  assign n5013 = n4897 & ~n5012;
  assign n5014 = ~n5006 & ~n5013;
  assign n5015 = ~n4712 & ~n4731;
  assign n5016 = ~n4722 & ~n4732;
  assign n5017 = ~n5015 & n5016;
  assign n5018 = ~n4721 & ~n5017;
  assign n5019 = ~n4736 & n5018;
  assign n5020 = n4937 & ~n5019;
  assign n5021 = ~n5014 & ~n5020;
  assign n5022 = ~n4980 & ~n5021;
  assign n5023 = pi00 & ~n4669;
  assign n5024 = ~pi01 & n5023;
  assign n5025 = ~n4961 & ~n4963;
  assign n5026 = ~n4946 & ~n4954;
  assign n5027 = ~n4953 & ~n4962;
  assign n5028 = ~pi02 & n4972;
  assign n5029 = ~n4973 & ~n5028;
  assign n5030 = n5025 & n5026;
  assign n5031 = n5027 & n5029;
  assign n5032 = n5030 & n5031;
  assign n5033 = n4939 & n5032;
  assign n5034 = ~n5024 & n5033;
  assign n5035 = ~n5022 & ~n5034;
  assign n5036 = n84 & n5033;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = n4698 & n5037;
  assign n5039 = ~n84 & ~n5024;
  assign n5040 = ~n4973 & ~n5039;
  assign n5041 = ~n5028 & ~n5040;
  assign n5042 = ~n4963 & n5041;
  assign n5043 = ~n4961 & ~n5042;
  assign n5044 = ~n4953 & ~n5043;
  assign n5045 = ~n4962 & ~n5044;
  assign n5046 = ~n4954 & ~n5045;
  assign n5047 = ~n4946 & ~n5046;
  assign n5048 = ~n4724 & ~n5047;
  assign n5049 = ~n4705 & ~n5048;
  assign n5050 = ~n4712 & n5049;
  assign n5051 = ~n4713 & ~n5050;
  assign n5052 = ~n4731 & ~n5051;
  assign n5053 = ~n4732 & ~n5052;
  assign n5054 = ~n4721 & ~n5053;
  assign n5055 = ~n4722 & ~n5054;
  assign n5056 = ~n4931 & ~n5055;
  assign n5057 = ~n4932 & ~n5056;
  assign n5058 = ~n4923 & n5057;
  assign n5059 = ~n4922 & ~n5058;
  assign n5060 = ~n4914 & ~n5059;
  assign n5061 = ~n4913 & ~n5060;
  assign n5062 = ~n4905 & ~n5061;
  assign n5063 = ~n4904 & ~n5062;
  assign n5064 = ~n4737 & ~n4883;
  assign n5065 = ~n5063 & n5064;
  assign n5066 = n5063 & ~n5064;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = ~n5037 & n5067;
  assign n5069 = ~n5038 & ~n5068;
  assign n5070 = ~n4705 & ~n4724;
  assign n5071 = ~n5047 & ~n5070;
  assign n5072 = n5047 & n5070;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = ~n5037 & ~n5073;
  assign n5075 = ~n4704 & n5037;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = pi07 & ~n5076;
  assign n5078 = n4720 & n5037;
  assign n5079 = n4723 & ~n5053;
  assign n5080 = ~n4723 & n5053;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = ~n5037 & n5081;
  assign n5083 = ~n5078 & ~n5082;
  assign n5084 = pi10 & n5083;
  assign n5085 = ~pi10 & ~n5083;
  assign n5086 = ~n5084 & ~n5085;
  assign n5087 = n4711 & n5037;
  assign n5088 = n4714 & ~n5049;
  assign n5089 = ~n4714 & n5049;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = ~n5037 & n5090;
  assign n5092 = ~n5087 & ~n5091;
  assign n5093 = pi08 & ~n5092;
  assign n5094 = ~pi08 & n5092;
  assign n5095 = ~n5093 & ~n5094;
  assign n5096 = ~pi07 & n5076;
  assign n5097 = ~n4733 & ~n5051;
  assign n5098 = n4733 & n5051;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = ~n5037 & ~n5099;
  assign n5101 = n4730 & n5037;
  assign n5102 = ~n5100 & ~n5101;
  assign n5103 = pi09 & n5102;
  assign n5104 = ~pi09 & ~n5102;
  assign n5105 = ~n5103 & ~n5104;
  assign n5106 = n5086 & ~n5096;
  assign n5107 = n5095 & n5105;
  assign n5108 = n5106 & n5107;
  assign n5109 = ~n4760 & n5037;
  assign n5110 = ~n4883 & ~n5063;
  assign n5111 = ~n4737 & ~n5110;
  assign n5112 = ~n4890 & n5111;
  assign n5113 = ~n4891 & ~n5112;
  assign n5114 = ~n4880 & ~n5113;
  assign n5115 = ~n4881 & ~n5114;
  assign n5116 = ~n4871 & ~n5115;
  assign n5117 = ~n4872 & ~n5116;
  assign n5118 = ~n4840 & ~n5117;
  assign n5119 = ~n4841 & ~n5118;
  assign n5120 = ~n4849 & ~n5119;
  assign n5121 = ~n4850 & ~n5120;
  assign n5122 = ~n4858 & ~n5121;
  assign n5123 = ~n4859 & ~n5122;
  assign n5124 = ~n4831 & ~n5123;
  assign n5125 = ~n4832 & ~n5124;
  assign n5126 = ~n4761 & ~n4808;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = n5125 & n5126;
  assign n5129 = ~n5037 & ~n5127;
  assign n5130 = ~n5128 & n5129;
  assign n5131 = ~n5109 & ~n5130;
  assign n5132 = pi23 & ~n5131;
  assign n5133 = ~pi23 & n5131;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = ~n4795 & n5037;
  assign n5136 = ~n4761 & ~n5125;
  assign n5137 = ~n4808 & ~n5136;
  assign n5138 = ~n4815 & ~n5137;
  assign n5139 = ~n4816 & ~n5138;
  assign n5140 = ~n4772 & ~n5139;
  assign n5141 = ~n4773 & ~n5140;
  assign n5142 = ~n4783 & ~n5141;
  assign n5143 = ~n4784 & ~n5142;
  assign n5144 = ~n4805 & ~n5143;
  assign n5145 = ~n4806 & ~n5144;
  assign n5146 = ~n4798 & ~n5145;
  assign n5147 = n4798 & n5145;
  assign n5148 = ~n5037 & ~n5146;
  assign n5149 = ~n5147 & n5148;
  assign n5150 = ~n5135 & ~n5149;
  assign n5151 = pi28 & ~n5150;
  assign n5152 = ~pi28 & n5150;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = ~n4785 & ~n5141;
  assign n5155 = n4785 & n5141;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = ~n5037 & ~n5156;
  assign n5158 = ~n4782 & n5037;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = pi26 & n5159;
  assign n5161 = ~pi26 & ~n5159;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = ~n4807 & ~n5143;
  assign n5164 = n4807 & n5143;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = ~n5037 & ~n5165;
  assign n5167 = ~n4804 & n5037;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = pi27 & n5168;
  assign n5170 = ~pi27 & ~n5168;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = ~n4774 & ~n5139;
  assign n5173 = n4774 & n5139;
  assign n5174 = ~n5172 & ~n5173;
  assign n5175 = ~n5037 & ~n5174;
  assign n5176 = ~n4771 & n5037;
  assign n5177 = ~n5175 & ~n5176;
  assign n5178 = pi25 & n5177;
  assign n5179 = ~pi25 & ~n5177;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = ~n4814 & n5037;
  assign n5182 = n4817 & ~n5137;
  assign n5183 = ~n4817 & n5137;
  assign n5184 = ~n5037 & ~n5182;
  assign n5185 = ~n5183 & n5184;
  assign n5186 = ~n5181 & ~n5185;
  assign n5187 = pi24 & n5186;
  assign n5188 = ~pi24 & ~n5186;
  assign n5189 = ~n5187 & ~n5188;
  assign n5190 = n67 & n5189;
  assign n5191 = n5180 & n5190;
  assign n5192 = n5162 & n5191;
  assign n5193 = n5171 & n5192;
  assign n5194 = n5153 & n5193;
  assign n5195 = n5134 & n5194;
  assign n5196 = ~n4830 & n5037;
  assign n5197 = n4833 & ~n5123;
  assign n5198 = ~n4833 & n5123;
  assign n5199 = ~n5037 & ~n5197;
  assign n5200 = ~n5198 & n5199;
  assign n5201 = ~n5196 & ~n5200;
  assign n5202 = pi22 & n5201;
  assign n5203 = ~pi22 & ~n5201;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = n4848 & n5037;
  assign n5206 = n4851 & ~n5119;
  assign n5207 = ~n4851 & n5119;
  assign n5208 = ~n5037 & ~n5206;
  assign n5209 = ~n5207 & n5208;
  assign n5210 = ~n5205 & ~n5209;
  assign n5211 = pi20 & n5210;
  assign n5212 = ~pi20 & ~n5210;
  assign n5213 = ~n5211 & ~n5212;
  assign n5214 = ~n4839 & n5037;
  assign n5215 = n4842 & ~n5117;
  assign n5216 = ~n4842 & n5117;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5037 & n5217;
  assign n5219 = ~n5214 & ~n5218;
  assign n5220 = pi19 & n5219;
  assign n5221 = ~pi19 & ~n5219;
  assign n5222 = ~n5220 & ~n5221;
  assign n5223 = ~n4857 & n5037;
  assign n5224 = ~n4860 & ~n5121;
  assign n5225 = n4860 & n5121;
  assign n5226 = ~n5037 & ~n5224;
  assign n5227 = ~n5225 & n5226;
  assign n5228 = ~n5223 & ~n5227;
  assign n5229 = pi21 & ~n5228;
  assign n5230 = ~pi21 & n5228;
  assign n5231 = ~n5229 & ~n5230;
  assign n5232 = n5213 & n5222;
  assign n5233 = n5231 & n5232;
  assign n5234 = n5204 & n5233;
  assign n5235 = n5195 & n5234;
  assign n5236 = ~n4882 & ~n5113;
  assign n5237 = n4882 & n5113;
  assign n5238 = ~n5236 & ~n5237;
  assign n5239 = ~n5037 & ~n5238;
  assign n5240 = ~n4879 & n5037;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = pi17 & n5241;
  assign n5243 = ~pi17 & ~n5241;
  assign n5244 = ~n5242 & ~n5243;
  assign n5245 = ~n4873 & ~n5115;
  assign n5246 = n4873 & n5115;
  assign n5247 = ~n5245 & ~n5246;
  assign n5248 = ~n5037 & ~n5247;
  assign n5249 = ~n4870 & n5037;
  assign n5250 = ~n5248 & ~n5249;
  assign n5251 = pi18 & n5250;
  assign n5252 = ~pi18 & ~n5250;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = n4889 & n5037;
  assign n5255 = n4892 & ~n5111;
  assign n5256 = ~n4892 & n5111;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = ~n5037 & n5257;
  assign n5259 = ~n5254 & ~n5258;
  assign n5260 = pi16 & ~n5259;
  assign n5261 = ~pi16 & n5259;
  assign n5262 = ~n5260 & ~n5261;
  assign n5263 = pi15 & ~n5069;
  assign n5264 = ~pi15 & n5069;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = n5244 & n5253;
  assign n5267 = n5262 & n5265;
  assign n5268 = n5266 & n5267;
  assign n5269 = n5235 & n5268;
  assign n5270 = n4903 & n5037;
  assign n5271 = ~n4906 & ~n5061;
  assign n5272 = n4906 & n5061;
  assign n5273 = ~n5271 & ~n5272;
  assign n5274 = ~n5037 & n5273;
  assign n5275 = ~n5270 & ~n5274;
  assign n5276 = pi14 & n5275;
  assign n5277 = ~pi14 & ~n5275;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = ~n4912 & n5037;
  assign n5280 = n4915 & ~n5059;
  assign n5281 = ~n4915 & n5059;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = ~n5037 & n5282;
  assign n5284 = ~n5279 & ~n5283;
  assign n5285 = pi13 & ~n5284;
  assign n5286 = ~pi13 & n5284;
  assign n5287 = ~n5285 & ~n5286;
  assign n5288 = ~n4921 & n5037;
  assign n5289 = ~n4924 & ~n5057;
  assign n5290 = n4924 & n5057;
  assign n5291 = ~n5289 & ~n5290;
  assign n5292 = ~n5037 & n5291;
  assign n5293 = ~n5288 & ~n5292;
  assign n5294 = pi12 & ~n5293;
  assign n5295 = ~pi12 & n5293;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = ~n4930 & n5037;
  assign n5298 = n4933 & ~n5055;
  assign n5299 = ~n4933 & n5055;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = ~n5037 & n5300;
  assign n5302 = ~n5297 & ~n5301;
  assign n5303 = pi11 & n5302;
  assign n5304 = ~pi11 & ~n5302;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = n5278 & n5287;
  assign n5307 = n5296 & n5305;
  assign n5308 = n5306 & n5307;
  assign n5309 = n5269 & n5308;
  assign n5310 = ~n5077 & n5108;
  assign n5311 = n5309 & n5310;
  assign n5312 = ~n4945 & n5037;
  assign n5313 = n5026 & ~n5045;
  assign n5314 = ~n5026 & n5045;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~n5037 & n5315;
  assign n5317 = ~n5312 & ~n5316;
  assign n5318 = pi06 & ~n5317;
  assign n5319 = ~n4952 & n5037;
  assign n5320 = n5027 & ~n5043;
  assign n5321 = ~n5027 & n5043;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = ~n5037 & n5322;
  assign n5324 = ~n5319 & ~n5323;
  assign n5325 = ~pi05 & n5324;
  assign n5326 = ~pi06 & n5317;
  assign n5327 = ~n4960 & n5037;
  assign n5328 = ~n5025 & ~n5041;
  assign n5329 = n5025 & n5041;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = ~n5037 & n5330;
  assign n5332 = ~n5327 & ~n5331;
  assign n5333 = pi04 & ~n5332;
  assign n5334 = pi05 & ~n5324;
  assign n5335 = ~pi04 & n5332;
  assign n5336 = ~n5029 & ~n5039;
  assign n5337 = n5029 & n5039;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = ~n5037 & ~n5338;
  assign n5340 = n4972 & n5037;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = pi03 & n5341;
  assign n5343 = ~n5335 & n5342;
  assign n5344 = ~n5333 & ~n5334;
  assign n5345 = ~n5343 & n5344;
  assign n5346 = ~n5325 & ~n5326;
  assign n5347 = ~n5345 & n5346;
  assign n5348 = ~n5318 & ~n5347;
  assign n5349 = n5311 & n5348;
  assign n5350 = ~n5212 & n5220;
  assign n5351 = ~n5211 & ~n5350;
  assign n5352 = ~n5229 & n5351;
  assign n5353 = ~n5230 & ~n5352;
  assign n5354 = ~n5203 & n5353;
  assign n5355 = ~n5202 & ~n5354;
  assign n5356 = n5195 & n5355;
  assign n5357 = ~n5133 & n5194;
  assign n5358 = ~n5178 & ~n5187;
  assign n5359 = ~n5179 & ~n5358;
  assign n5360 = ~n5161 & n5359;
  assign n5361 = ~n5160 & ~n5360;
  assign n5362 = ~n5169 & n5361;
  assign n5363 = ~n5170 & ~n5362;
  assign n5364 = ~n5152 & n5363;
  assign n5365 = n67 & ~n5151;
  assign n5366 = ~n5364 & n5365;
  assign n5367 = ~n5357 & n5366;
  assign n5368 = ~n5356 & ~n5367;
  assign n5369 = ~n5261 & ~n5264;
  assign n5370 = ~n5242 & ~n5260;
  assign n5371 = ~n5369 & n5370;
  assign n5372 = ~n5243 & ~n5252;
  assign n5373 = ~n5371 & n5372;
  assign n5374 = ~n5251 & ~n5373;
  assign n5375 = n5235 & ~n5374;
  assign n5376 = ~n5368 & ~n5375;
  assign n5377 = ~n5294 & ~n5303;
  assign n5378 = ~n5286 & ~n5295;
  assign n5379 = ~n5377 & n5378;
  assign n5380 = ~n5276 & ~n5285;
  assign n5381 = ~n5379 & n5380;
  assign n5382 = ~n5277 & ~n5381;
  assign n5383 = n5269 & ~n5382;
  assign n5384 = ~n5376 & ~n5383;
  assign n5385 = n5093 & ~n5104;
  assign n5386 = ~n5084 & ~n5103;
  assign n5387 = ~n5385 & n5386;
  assign n5388 = ~n5085 & ~n5387;
  assign n5389 = ~n5108 & ~n5388;
  assign n5390 = n5309 & ~n5389;
  assign n5391 = ~n5384 & ~n5390;
  assign n5392 = ~n5349 & ~n5391;
  assign n5393 = n314 & n4661;
  assign n5394 = pi01 & ~n4661;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~n5037 & n5395;
  assign n5397 = ~n5023 & n5037;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = pi02 & ~n5398;
  assign n5400 = ~pi02 & n5398;
  assign n5401 = pi00 & n5035;
  assign n5402 = ~pi01 & n5401;
  assign n5403 = ~n5400 & ~n5402;
  assign n5404 = ~n5399 & ~n5403;
  assign n5405 = ~n5333 & ~n5335;
  assign n5406 = ~n5318 & ~n5326;
  assign n5407 = ~n5325 & ~n5334;
  assign n5408 = ~pi03 & ~n5341;
  assign n5409 = ~n5342 & ~n5408;
  assign n5410 = n5405 & n5406;
  assign n5411 = n5407 & n5409;
  assign n5412 = n5410 & n5411;
  assign n5413 = n5311 & n5412;
  assign n5414 = ~n5404 & n5413;
  assign n5415 = ~n5392 & ~n5414;
  assign n5416 = ~n5399 & ~n5400;
  assign n5417 = n84 & n5416;
  assign n5418 = n5413 & n5417;
  assign n5419 = ~n5415 & ~n5418;
  assign n5420 = n5069 & n5419;
  assign n5421 = pi00 & ~n5035;
  assign n5422 = ~pi01 & ~n5421;
  assign n5423 = ~n5400 & ~n5422;
  assign n5424 = ~n5399 & ~n5423;
  assign n5425 = ~n5342 & n5424;
  assign n5426 = ~n5408 & ~n5425;
  assign n5427 = ~n5335 & n5426;
  assign n5428 = ~n5333 & ~n5427;
  assign n5429 = ~n5325 & ~n5428;
  assign n5430 = ~n5334 & ~n5429;
  assign n5431 = ~n5326 & ~n5430;
  assign n5432 = ~n5318 & ~n5431;
  assign n5433 = ~n5096 & ~n5432;
  assign n5434 = ~n5077 & ~n5433;
  assign n5435 = ~n5094 & ~n5434;
  assign n5436 = ~n5093 & ~n5435;
  assign n5437 = ~n5104 & ~n5436;
  assign n5438 = ~n5103 & ~n5437;
  assign n5439 = ~n5084 & n5438;
  assign n5440 = ~n5085 & ~n5439;
  assign n5441 = ~n5303 & ~n5440;
  assign n5442 = ~n5304 & ~n5441;
  assign n5443 = ~n5295 & n5442;
  assign n5444 = ~n5294 & ~n5443;
  assign n5445 = ~n5286 & ~n5444;
  assign n5446 = ~n5285 & ~n5445;
  assign n5447 = ~n5276 & n5446;
  assign n5448 = ~n5277 & ~n5447;
  assign n5449 = n5265 & ~n5448;
  assign n5450 = ~n5265 & n5448;
  assign n5451 = ~n5449 & ~n5450;
  assign n5452 = ~n5419 & n5451;
  assign n5453 = ~n5420 & ~n5452;
  assign n5454 = n5250 & n5419;
  assign n5455 = ~n5264 & n5448;
  assign n5456 = ~n5263 & ~n5455;
  assign n5457 = ~n5261 & ~n5456;
  assign n5458 = ~n5260 & ~n5457;
  assign n5459 = ~n5243 & ~n5458;
  assign n5460 = ~n5242 & ~n5459;
  assign n5461 = n5253 & ~n5460;
  assign n5462 = ~n5253 & n5460;
  assign n5463 = ~n5419 & ~n5461;
  assign n5464 = ~n5462 & n5463;
  assign n5465 = ~n5454 & ~n5464;
  assign n5466 = ~pi19 & n5465;
  assign n5467 = pi19 & ~n5465;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = n5131 & n5419;
  assign n5470 = ~n5252 & ~n5460;
  assign n5471 = ~n5251 & ~n5470;
  assign n5472 = ~n5220 & n5471;
  assign n5473 = ~n5221 & ~n5472;
  assign n5474 = ~n5211 & ~n5473;
  assign n5475 = ~n5212 & ~n5474;
  assign n5476 = ~n5229 & ~n5475;
  assign n5477 = ~n5230 & ~n5476;
  assign n5478 = ~n5202 & ~n5477;
  assign n5479 = ~n5203 & ~n5478;
  assign n5480 = n5134 & ~n5479;
  assign n5481 = ~n5134 & n5479;
  assign n5482 = ~n5419 & ~n5480;
  assign n5483 = ~n5481 & n5482;
  assign n5484 = ~n5469 & ~n5483;
  assign n5485 = pi24 & n5484;
  assign n5486 = ~n5150 & n5419;
  assign n5487 = ~n5133 & n5479;
  assign n5488 = ~n5132 & ~n5487;
  assign n5489 = ~n5188 & ~n5488;
  assign n5490 = ~n5187 & ~n5489;
  assign n5491 = ~n5178 & n5490;
  assign n5492 = ~n5179 & ~n5491;
  assign n5493 = ~n5160 & ~n5492;
  assign n5494 = ~n5161 & ~n5493;
  assign n5495 = ~n5169 & ~n5494;
  assign n5496 = ~n5170 & ~n5495;
  assign n5497 = ~n5153 & ~n5496;
  assign n5498 = n5153 & n5496;
  assign n5499 = ~n5419 & ~n5497;
  assign n5500 = ~n5498 & n5499;
  assign n5501 = ~n5486 & ~n5500;
  assign n5502 = ~pi29 & n5501;
  assign n5503 = pi29 & ~n5501;
  assign n5504 = ~n5502 & ~n5503;
  assign n5505 = ~n5171 & ~n5494;
  assign n5506 = n5171 & n5494;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = ~n5419 & ~n5507;
  assign n5509 = ~n5168 & n5419;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = pi28 & n5510;
  assign n5512 = ~pi28 & ~n5510;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = n5177 & n5419;
  assign n5515 = n5180 & ~n5490;
  assign n5516 = ~n5180 & n5490;
  assign n5517 = ~n5419 & ~n5515;
  assign n5518 = ~n5516 & n5517;
  assign n5519 = ~n5514 & ~n5518;
  assign n5520 = ~pi26 & n5519;
  assign n5521 = pi26 & ~n5519;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = ~n5189 & ~n5488;
  assign n5524 = n5189 & n5488;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = ~n5419 & ~n5525;
  assign n5527 = n5186 & n5419;
  assign n5528 = ~n5526 & ~n5527;
  assign n5529 = pi25 & ~n5528;
  assign n5530 = ~pi25 & n5528;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = ~pi24 & ~n5484;
  assign n5533 = ~n5162 & ~n5492;
  assign n5534 = n5162 & n5492;
  assign n5535 = ~n5533 & ~n5534;
  assign n5536 = ~n5419 & ~n5535;
  assign n5537 = ~n5159 & n5419;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = pi27 & n5538;
  assign n5540 = ~pi27 & ~n5538;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = n66 & ~n5532;
  assign n5543 = n5531 & n5542;
  assign n5544 = n5522 & n5543;
  assign n5545 = n5541 & n5544;
  assign n5546 = n5513 & n5545;
  assign n5547 = n5504 & n5546;
  assign n5548 = ~n5485 & n5547;
  assign n5549 = ~n5204 & ~n5477;
  assign n5550 = n5204 & n5477;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = ~n5419 & ~n5551;
  assign n5553 = ~n5201 & n5419;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = pi23 & n5554;
  assign n5556 = ~pi23 & ~n5554;
  assign n5557 = ~n5555 & ~n5556;
  assign n5558 = ~n5210 & n5419;
  assign n5559 = n5213 & ~n5473;
  assign n5560 = ~n5213 & n5473;
  assign n5561 = ~n5419 & ~n5559;
  assign n5562 = ~n5560 & n5561;
  assign n5563 = ~n5558 & ~n5562;
  assign n5564 = pi21 & n5563;
  assign n5565 = ~pi21 & ~n5563;
  assign n5566 = ~n5564 & ~n5565;
  assign n5567 = n5219 & n5419;
  assign n5568 = n5222 & ~n5471;
  assign n5569 = ~n5222 & n5471;
  assign n5570 = ~n5419 & ~n5568;
  assign n5571 = ~n5569 & n5570;
  assign n5572 = ~n5567 & ~n5571;
  assign n5573 = pi20 & ~n5572;
  assign n5574 = ~pi20 & n5572;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 = n5228 & n5419;
  assign n5577 = n5231 & ~n5475;
  assign n5578 = ~n5231 & n5475;
  assign n5579 = ~n5419 & ~n5577;
  assign n5580 = ~n5578 & n5579;
  assign n5581 = ~n5576 & ~n5580;
  assign n5582 = ~pi22 & ~n5581;
  assign n5583 = pi22 & n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = n5566 & n5575;
  assign n5586 = n5584 & n5585;
  assign n5587 = n5557 & n5586;
  assign n5588 = n5548 & n5587;
  assign n5589 = ~pi16 & ~n5453;
  assign n5590 = pi16 & n5453;
  assign n5591 = ~n5589 & ~n5590;
  assign n5592 = n5241 & n5419;
  assign n5593 = n5244 & ~n5458;
  assign n5594 = ~n5244 & n5458;
  assign n5595 = ~n5419 & ~n5593;
  assign n5596 = ~n5594 & n5595;
  assign n5597 = ~n5592 & ~n5596;
  assign n5598 = pi18 & ~n5597;
  assign n5599 = ~pi18 & n5597;
  assign n5600 = ~n5598 & ~n5599;
  assign n5601 = ~n5262 & ~n5456;
  assign n5602 = n5262 & n5456;
  assign n5603 = ~n5601 & ~n5602;
  assign n5604 = ~n5419 & ~n5603;
  assign n5605 = ~n5259 & n5419;
  assign n5606 = ~n5604 & ~n5605;
  assign n5607 = ~pi17 & n5606;
  assign n5608 = pi17 & ~n5606;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = n5591 & n5609;
  assign n5611 = n5600 & n5610;
  assign n5612 = n5468 & n5611;
  assign n5613 = n5588 & n5612;
  assign n5614 = n5275 & n5419;
  assign n5615 = n5278 & ~n5446;
  assign n5616 = ~n5278 & n5446;
  assign n5617 = ~n5615 & ~n5616;
  assign n5618 = ~n5419 & n5617;
  assign n5619 = ~n5614 & ~n5618;
  assign n5620 = pi15 & ~n5619;
  assign n5621 = ~pi15 & n5619;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = ~n5284 & n5419;
  assign n5624 = n5287 & ~n5444;
  assign n5625 = ~n5287 & n5444;
  assign n5626 = ~n5624 & ~n5625;
  assign n5627 = ~n5419 & n5626;
  assign n5628 = ~n5623 & ~n5627;
  assign n5629 = pi14 & ~n5628;
  assign n5630 = ~pi14 & n5628;
  assign n5631 = ~n5629 & ~n5630;
  assign n5632 = n5293 & n5419;
  assign n5633 = n5296 & ~n5442;
  assign n5634 = ~n5296 & n5442;
  assign n5635 = ~n5633 & ~n5634;
  assign n5636 = ~n5419 & n5635;
  assign n5637 = ~n5632 & ~n5636;
  assign n5638 = pi13 & n5637;
  assign n5639 = ~pi13 & ~n5637;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = ~n5302 & n5419;
  assign n5642 = n5305 & ~n5440;
  assign n5643 = ~n5305 & n5440;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = ~n5419 & n5644;
  assign n5646 = ~n5641 & ~n5645;
  assign n5647 = pi12 & n5646;
  assign n5648 = ~pi12 & ~n5646;
  assign n5649 = ~n5647 & ~n5648;
  assign n5650 = n5622 & n5631;
  assign n5651 = n5640 & n5649;
  assign n5652 = n5650 & n5651;
  assign n5653 = n5613 & n5652;
  assign n5654 = n5083 & n5419;
  assign n5655 = n5086 & ~n5438;
  assign n5656 = ~n5086 & n5438;
  assign n5657 = ~n5655 & ~n5656;
  assign n5658 = ~n5419 & n5657;
  assign n5659 = ~n5654 & ~n5658;
  assign n5660 = ~pi11 & n5659;
  assign n5661 = pi11 & ~n5659;
  assign n5662 = n5102 & n5419;
  assign n5663 = n5105 & ~n5436;
  assign n5664 = ~n5105 & n5436;
  assign n5665 = ~n5663 & ~n5664;
  assign n5666 = ~n5419 & n5665;
  assign n5667 = ~n5662 & ~n5666;
  assign n5668 = pi10 & ~n5667;
  assign n5669 = ~n5092 & n5419;
  assign n5670 = n5095 & ~n5434;
  assign n5671 = ~n5095 & n5434;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = ~n5419 & n5672;
  assign n5674 = ~n5669 & ~n5673;
  assign n5675 = ~pi09 & n5674;
  assign n5676 = ~pi10 & n5667;
  assign n5677 = ~n5077 & ~n5096;
  assign n5678 = ~n5432 & ~n5677;
  assign n5679 = n5432 & n5677;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = ~n5419 & ~n5680;
  assign n5682 = ~n5076 & n5419;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = ~pi08 & n5683;
  assign n5685 = pi09 & ~n5674;
  assign n5686 = n5684 & ~n5685;
  assign n5687 = ~n5675 & ~n5676;
  assign n5688 = ~n5686 & n5687;
  assign n5689 = ~n5661 & ~n5668;
  assign n5690 = ~n5688 & n5689;
  assign n5691 = ~n5660 & ~n5690;
  assign n5692 = n5653 & n5691;
  assign n5693 = ~n5638 & ~n5647;
  assign n5694 = ~n5630 & ~n5639;
  assign n5695 = ~n5693 & n5694;
  assign n5696 = ~n5620 & ~n5629;
  assign n5697 = ~n5695 & n5696;
  assign n5698 = ~n5621 & ~n5697;
  assign n5699 = n5613 & ~n5698;
  assign n5700 = ~n5520 & n5529;
  assign n5701 = ~n5521 & ~n5700;
  assign n5702 = ~n5539 & n5701;
  assign n5703 = ~n5540 & ~n5702;
  assign n5704 = ~n5512 & n5703;
  assign n5705 = ~n5511 & ~n5704;
  assign n5706 = ~n5502 & ~n5705;
  assign n5707 = n66 & ~n5503;
  assign n5708 = ~n5706 & n5707;
  assign n5709 = ~n5547 & n5708;
  assign n5710 = ~n5565 & n5573;
  assign n5711 = ~n5564 & ~n5710;
  assign n5712 = ~n5583 & n5711;
  assign n5713 = ~n5582 & ~n5712;
  assign n5714 = ~n5556 & n5713;
  assign n5715 = ~n5555 & ~n5714;
  assign n5716 = n5548 & n5715;
  assign n5717 = ~n5588 & ~n5709;
  assign n5718 = ~n5716 & n5717;
  assign n5719 = n5589 & ~n5608;
  assign n5720 = ~n5607 & ~n5719;
  assign n5721 = ~n5599 & n5720;
  assign n5722 = ~n5598 & ~n5721;
  assign n5723 = ~n5467 & n5722;
  assign n5724 = ~n5466 & ~n5723;
  assign n5725 = n5588 & n5724;
  assign n5726 = ~n5718 & ~n5725;
  assign n5727 = ~n5699 & ~n5726;
  assign n5728 = ~n5692 & ~n5727;
  assign n5729 = ~n5660 & ~n5661;
  assign n5730 = pi08 & ~n5683;
  assign n5731 = ~n5684 & ~n5730;
  assign n5732 = ~n5675 & ~n5685;
  assign n5733 = ~n5668 & ~n5676;
  assign n5734 = n5729 & n5731;
  assign n5735 = n5732 & n5733;
  assign n5736 = n5734 & n5735;
  assign n5737 = n5653 & n5736;
  assign n5738 = ~n5317 & n5419;
  assign n5739 = n5406 & ~n5430;
  assign n5740 = ~n5406 & n5430;
  assign n5741 = ~n5739 & ~n5740;
  assign n5742 = ~n5419 & n5741;
  assign n5743 = ~n5738 & ~n5742;
  assign n5744 = ~pi07 & n5743;
  assign n5745 = pi07 & ~n5743;
  assign n5746 = ~n5324 & n5419;
  assign n5747 = n5407 & ~n5428;
  assign n5748 = ~n5407 & n5428;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = ~n5419 & n5749;
  assign n5751 = ~n5746 & ~n5750;
  assign n5752 = ~pi06 & n5751;
  assign n5753 = ~n5332 & n5419;
  assign n5754 = ~n5405 & ~n5426;
  assign n5755 = n5405 & n5426;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = ~n5419 & n5756;
  assign n5758 = ~n5753 & ~n5757;
  assign n5759 = pi05 & ~n5758;
  assign n5760 = pi06 & ~n5751;
  assign n5761 = n5341 & n5419;
  assign n5762 = n5409 & ~n5424;
  assign n5763 = ~n5409 & n5424;
  assign n5764 = ~n5762 & ~n5763;
  assign n5765 = ~n5419 & n5764;
  assign n5766 = ~n5761 & ~n5765;
  assign n5767 = pi04 & ~n5766;
  assign n5768 = ~pi05 & n5758;
  assign n5769 = n5767 & ~n5768;
  assign n5770 = ~n5759 & ~n5760;
  assign n5771 = ~n5769 & n5770;
  assign n5772 = ~n5752 & ~n5771;
  assign n5773 = ~n5745 & ~n5772;
  assign n5774 = ~n5744 & ~n5773;
  assign n5775 = n5737 & ~n5774;
  assign n5776 = ~n5728 & ~n5775;
  assign n5777 = ~n5752 & ~n5760;
  assign n5778 = ~n5759 & ~n5768;
  assign n5779 = ~n5744 & ~n5745;
  assign n5780 = ~pi04 & n5766;
  assign n5781 = ~n5767 & ~n5780;
  assign n5782 = n5777 & n5778;
  assign n5783 = n5779 & n5781;
  assign n5784 = n5782 & n5783;
  assign n5785 = n5737 & n5784;
  assign n5786 = n5398 & n5419;
  assign n5787 = ~n5416 & ~n5422;
  assign n5788 = n5416 & n5422;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = ~n5419 & n5789;
  assign n5791 = ~n5786 & ~n5790;
  assign n5792 = pi03 & n5791;
  assign n5793 = n314 & ~n5419;
  assign n5794 = ~n5401 & ~n5793;
  assign n5795 = n5402 & ~n5419;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = ~pi02 & n5796;
  assign n5798 = pi02 & ~n5796;
  assign n5799 = pi00 & ~n5419;
  assign n5800 = ~pi01 & n5799;
  assign n5801 = ~n5798 & n5800;
  assign n5802 = ~pi03 & ~n5791;
  assign n5803 = ~n5797 & ~n5802;
  assign n5804 = ~n5801 & n5803;
  assign n5805 = ~n5792 & ~n5804;
  assign n5806 = n5785 & ~n5805;
  assign n5807 = ~n5776 & ~n5806;
  assign n5808 = ~n5797 & ~n5798;
  assign n5809 = ~n5792 & ~n5802;
  assign n5810 = n84 & n5809;
  assign n5811 = n5808 & n5810;
  assign n5812 = n5785 & n5811;
  assign n5813 = ~n5807 & ~n5812;
  assign n5814 = n5453 & n5813;
  assign n5815 = ~n84 & ~n5800;
  assign n5816 = ~n5797 & n5815;
  assign n5817 = ~n5798 & ~n5816;
  assign n5818 = ~n5802 & ~n5817;
  assign n5819 = ~n5792 & ~n5818;
  assign n5820 = ~n5780 & ~n5819;
  assign n5821 = ~n5767 & ~n5820;
  assign n5822 = ~n5768 & ~n5821;
  assign n5823 = ~n5759 & ~n5822;
  assign n5824 = ~n5752 & ~n5823;
  assign n5825 = ~n5760 & ~n5824;
  assign n5826 = ~n5744 & ~n5825;
  assign n5827 = ~n5745 & ~n5826;
  assign n5828 = ~n5684 & ~n5827;
  assign n5829 = ~n5730 & ~n5828;
  assign n5830 = ~n5675 & ~n5829;
  assign n5831 = ~n5685 & ~n5830;
  assign n5832 = ~n5676 & ~n5831;
  assign n5833 = ~n5668 & ~n5832;
  assign n5834 = ~n5660 & ~n5833;
  assign n5835 = ~n5661 & ~n5834;
  assign n5836 = ~n5648 & ~n5835;
  assign n5837 = ~n5647 & ~n5836;
  assign n5838 = ~n5638 & n5837;
  assign n5839 = ~n5639 & ~n5838;
  assign n5840 = ~n5630 & n5839;
  assign n5841 = ~n5629 & ~n5840;
  assign n5842 = ~n5621 & ~n5841;
  assign n5843 = ~n5620 & ~n5842;
  assign n5844 = n5591 & ~n5843;
  assign n5845 = ~n5591 & n5843;
  assign n5846 = ~n5844 & ~n5845;
  assign n5847 = ~n5813 & n5846;
  assign n5848 = ~n5814 & ~n5847;
  assign n5849 = ~n5796 & n5813;
  assign n5850 = ~n5808 & ~n5815;
  assign n5851 = n5808 & n5815;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n5813 & n5852;
  assign n5854 = ~n5849 & ~n5853;
  assign n5855 = pi03 & ~n5854;
  assign n5856 = ~pi03 & n5854;
  assign n5857 = ~n5855 & ~n5856;
  assign n5858 = n5791 & n5813;
  assign n5859 = n5809 & ~n5817;
  assign n5860 = ~n5809 & n5817;
  assign n5861 = ~n5859 & ~n5860;
  assign n5862 = ~n5813 & n5861;
  assign n5863 = ~n5858 & ~n5862;
  assign n5864 = pi04 & ~n5863;
  assign n5865 = ~pi04 & n5863;
  assign n5866 = ~n5864 & ~n5865;
  assign n5867 = n5538 & n5813;
  assign n5868 = ~n5589 & ~n5843;
  assign n5869 = ~n5590 & ~n5868;
  assign n5870 = ~n5607 & ~n5869;
  assign n5871 = ~n5608 & ~n5870;
  assign n5872 = ~n5599 & ~n5871;
  assign n5873 = ~n5598 & ~n5872;
  assign n5874 = ~n5466 & ~n5873;
  assign n5875 = ~n5467 & ~n5874;
  assign n5876 = ~n5574 & ~n5875;
  assign n5877 = ~n5573 & ~n5876;
  assign n5878 = ~n5565 & ~n5877;
  assign n5879 = ~n5564 & ~n5878;
  assign n5880 = ~n5583 & n5879;
  assign n5881 = ~n5582 & ~n5880;
  assign n5882 = ~n5555 & ~n5881;
  assign n5883 = ~n5556 & ~n5882;
  assign n5884 = ~n5485 & ~n5883;
  assign n5885 = ~n5532 & ~n5884;
  assign n5886 = ~n5530 & n5885;
  assign n5887 = ~n5529 & ~n5886;
  assign n5888 = ~n5520 & ~n5887;
  assign n5889 = ~n5521 & ~n5888;
  assign n5890 = n5541 & ~n5889;
  assign n5891 = ~n5541 & n5889;
  assign n5892 = ~n5813 & ~n5890;
  assign n5893 = ~n5891 & n5892;
  assign n5894 = ~n5867 & ~n5893;
  assign n5895 = ~pi28 & n5894;
  assign n5896 = pi28 & ~n5894;
  assign n5897 = ~n5895 & ~n5896;
  assign n5898 = n5519 & n5813;
  assign n5899 = ~n5522 & ~n5887;
  assign n5900 = n5522 & n5887;
  assign n5901 = ~n5813 & ~n5899;
  assign n5902 = ~n5900 & n5901;
  assign n5903 = ~n5898 & ~n5902;
  assign n5904 = ~pi27 & ~n5903;
  assign n5905 = pi27 & n5903;
  assign n5906 = ~n5904 & ~n5905;
  assign n5907 = ~n5484 & n5813;
  assign n5908 = ~n5485 & ~n5532;
  assign n5909 = n5883 & ~n5908;
  assign n5910 = ~n5883 & n5908;
  assign n5911 = ~n5813 & ~n5909;
  assign n5912 = ~n5910 & n5911;
  assign n5913 = ~n5907 & ~n5912;
  assign n5914 = ~pi25 & ~n5913;
  assign n5915 = ~n5528 & n5813;
  assign n5916 = ~n5531 & ~n5885;
  assign n5917 = n5531 & n5885;
  assign n5918 = ~n5813 & ~n5916;
  assign n5919 = ~n5917 & n5918;
  assign n5920 = ~n5915 & ~n5919;
  assign n5921 = pi26 & ~n5920;
  assign n5922 = ~pi26 & n5920;
  assign n5923 = ~n5921 & ~n5922;
  assign n5924 = ~pi31 & ~n5914;
  assign n5925 = n5923 & n5924;
  assign n5926 = n5906 & n5925;
  assign n5927 = ~n5501 & n5813;
  assign n5928 = ~n5539 & n5889;
  assign n5929 = ~n5540 & ~n5928;
  assign n5930 = ~n5511 & ~n5929;
  assign n5931 = ~n5512 & ~n5930;
  assign n5932 = ~n5504 & ~n5931;
  assign n5933 = n5504 & n5931;
  assign n5934 = ~n5813 & ~n5932;
  assign n5935 = ~n5933 & n5934;
  assign n5936 = ~n5927 & ~n5935;
  assign n5937 = ~pi30 & n5936;
  assign n5938 = pi30 & ~n5936;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = ~n5513 & ~n5929;
  assign n5941 = n5513 & n5929;
  assign n5942 = ~n5940 & ~n5941;
  assign n5943 = ~n5813 & ~n5942;
  assign n5944 = ~n5510 & n5813;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = pi29 & n5945;
  assign n5947 = ~pi29 & ~n5945;
  assign n5948 = ~n5946 & ~n5947;
  assign n5949 = pi25 & n5913;
  assign n5950 = n5926 & ~n5949;
  assign n5951 = n5897 & n5950;
  assign n5952 = n5948 & n5951;
  assign n5953 = n5939 & n5952;
  assign n5954 = ~n5554 & n5813;
  assign n5955 = n5557 & ~n5881;
  assign n5956 = ~n5557 & n5881;
  assign n5957 = ~n5813 & ~n5955;
  assign n5958 = ~n5956 & n5957;
  assign n5959 = ~n5954 & ~n5958;
  assign n5960 = pi24 & n5959;
  assign n5961 = ~pi24 & ~n5959;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n5572 & n5813;
  assign n5964 = n5575 & ~n5875;
  assign n5965 = ~n5575 & n5875;
  assign n5966 = ~n5813 & ~n5964;
  assign n5967 = ~n5965 & n5966;
  assign n5968 = ~n5963 & ~n5967;
  assign n5969 = pi21 & ~n5968;
  assign n5970 = ~pi21 & n5968;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = n5563 & n5813;
  assign n5973 = n5566 & ~n5877;
  assign n5974 = ~n5566 & n5877;
  assign n5975 = ~n5813 & ~n5973;
  assign n5976 = ~n5974 & n5975;
  assign n5977 = ~n5972 & ~n5976;
  assign n5978 = pi22 & ~n5977;
  assign n5979 = ~pi22 & n5977;
  assign n5980 = ~n5978 & ~n5979;
  assign n5981 = ~n5584 & ~n5879;
  assign n5982 = n5584 & n5879;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5813 & ~n5983;
  assign n5985 = n5581 & n5813;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = ~pi23 & n5986;
  assign n5988 = pi23 & ~n5986;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = n5971 & n5980;
  assign n5991 = n5989 & n5990;
  assign n5992 = n5962 & n5991;
  assign n5993 = n5953 & n5992;
  assign n5994 = ~n5465 & n5813;
  assign n5995 = n5468 & ~n5873;
  assign n5996 = ~n5468 & n5873;
  assign n5997 = ~n5995 & ~n5996;
  assign n5998 = ~n5813 & n5997;
  assign n5999 = ~n5994 & ~n5998;
  assign n6000 = ~pi20 & n5999;
  assign n6001 = pi20 & ~n5999;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n5606 & n5813;
  assign n6004 = n5609 & ~n5869;
  assign n6005 = ~n5609 & n5869;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = ~n5813 & n6006;
  assign n6008 = ~n6003 & ~n6007;
  assign n6009 = ~pi18 & n6008;
  assign n6010 = pi18 & ~n6008;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = ~n5600 & ~n5871;
  assign n6013 = n5600 & n5871;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = ~n5813 & ~n6014;
  assign n6016 = ~n5597 & n5813;
  assign n6017 = ~n6015 & ~n6016;
  assign n6018 = pi19 & ~n6017;
  assign n6019 = ~pi19 & n6017;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = ~pi17 & n5848;
  assign n6022 = pi17 & ~n5848;
  assign n6023 = ~n6021 & ~n6022;
  assign n6024 = n6002 & n6011;
  assign n6025 = n6020 & n6023;
  assign n6026 = n6024 & n6025;
  assign n6027 = n5993 & n6026;
  assign n6028 = n5619 & n5813;
  assign n6029 = ~n5622 & ~n5841;
  assign n6030 = n5622 & n5841;
  assign n6031 = ~n6029 & ~n6030;
  assign n6032 = ~n5813 & n6031;
  assign n6033 = ~n6028 & ~n6032;
  assign n6034 = pi16 & n6033;
  assign n6035 = ~pi16 & ~n6033;
  assign n6036 = ~n6034 & ~n6035;
  assign n6037 = ~n5628 & n5813;
  assign n6038 = ~n5631 & ~n5839;
  assign n6039 = n5631 & n5839;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = ~n5813 & n6040;
  assign n6042 = ~n6037 & ~n6041;
  assign n6043 = ~pi15 & n6042;
  assign n6044 = pi15 & ~n6042;
  assign n6045 = ~n6043 & ~n6044;
  assign n6046 = ~n5640 & ~n5837;
  assign n6047 = n5640 & n5837;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = ~n5813 & ~n6048;
  assign n6050 = n5637 & n5813;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = pi14 & ~n6051;
  assign n6053 = ~pi14 & n6051;
  assign n6054 = ~n6052 & ~n6053;
  assign n6055 = n5646 & n5813;
  assign n6056 = n5649 & ~n5835;
  assign n6057 = ~n5649 & n5835;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = ~n5813 & n6058;
  assign n6060 = ~n6055 & ~n6059;
  assign n6061 = pi13 & ~n6060;
  assign n6062 = ~pi13 & n6060;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = n6036 & n6045;
  assign n6065 = n6054 & n6063;
  assign n6066 = n6064 & n6065;
  assign n6067 = n6027 & n6066;
  assign n6068 = ~n5667 & n5813;
  assign n6069 = n5733 & ~n5831;
  assign n6070 = ~n5733 & n5831;
  assign n6071 = ~n6069 & ~n6070;
  assign n6072 = ~n5813 & n6071;
  assign n6073 = ~n6068 & ~n6072;
  assign n6074 = pi11 & ~n6073;
  assign n6075 = ~pi11 & n6073;
  assign n6076 = ~n6074 & ~n6075;
  assign n6077 = ~n5674 & n5813;
  assign n6078 = n5732 & ~n5829;
  assign n6079 = ~n5732 & n5829;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = ~n5813 & n6080;
  assign n6082 = ~n6077 & ~n6081;
  assign n6083 = pi10 & ~n6082;
  assign n6084 = ~pi10 & n6082;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = ~n5683 & n5813;
  assign n6087 = n5731 & ~n5827;
  assign n6088 = ~n5731 & n5827;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = ~n5813 & n6089;
  assign n6091 = ~n6086 & ~n6090;
  assign n6092 = ~pi09 & n6091;
  assign n6093 = pi09 & ~n6091;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = ~n5659 & n5813;
  assign n6096 = n5729 & ~n5833;
  assign n6097 = ~n5729 & n5833;
  assign n6098 = ~n6096 & ~n6097;
  assign n6099 = ~n5813 & n6098;
  assign n6100 = ~n6095 & ~n6099;
  assign n6101 = ~pi12 & n6100;
  assign n6102 = pi12 & ~n6100;
  assign n6103 = ~n6101 & ~n6102;
  assign n6104 = n6076 & n6085;
  assign n6105 = n6094 & n6103;
  assign n6106 = n6104 & n6105;
  assign n6107 = n6067 & n6106;
  assign n6108 = ~n5743 & n5813;
  assign n6109 = n5779 & ~n5825;
  assign n6110 = ~n5779 & n5825;
  assign n6111 = ~n6109 & ~n6110;
  assign n6112 = ~n5813 & n6111;
  assign n6113 = ~n6108 & ~n6112;
  assign n6114 = pi08 & ~n6113;
  assign n6115 = ~pi08 & n6113;
  assign n6116 = ~n6114 & ~n6115;
  assign n6117 = ~n5751 & n5813;
  assign n6118 = n5777 & ~n5823;
  assign n6119 = ~n5777 & n5823;
  assign n6120 = ~n6118 & ~n6119;
  assign n6121 = ~n5813 & n6120;
  assign n6122 = ~n6117 & ~n6121;
  assign n6123 = pi07 & ~n6122;
  assign n6124 = ~pi07 & n6122;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = ~n5758 & n5813;
  assign n6127 = n5778 & ~n5821;
  assign n6128 = ~n5778 & n5821;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = ~n5813 & n6129;
  assign n6131 = ~n6126 & ~n6130;
  assign n6132 = ~pi06 & n6131;
  assign n6133 = pi06 & ~n6131;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = ~n5766 & n5813;
  assign n6136 = n5781 & ~n5819;
  assign n6137 = ~n5781 & n5819;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = ~n5813 & n6138;
  assign n6140 = ~n6135 & ~n6139;
  assign n6141 = pi05 & ~n6140;
  assign n6142 = ~pi05 & n6140;
  assign n6143 = ~n6141 & ~n6142;
  assign n6144 = n6116 & n6125;
  assign n6145 = n6134 & n6143;
  assign n6146 = n6144 & n6145;
  assign n6147 = n6107 & n6146;
  assign n6148 = n5857 & n5866;
  assign n6149 = n6147 & n6148;
  assign n6150 = pi00 & ~n5415;
  assign n6151 = ~pi01 & ~n6150;
  assign n6152 = pi01 & n6150;
  assign n6153 = ~n6151 & ~n6152;
  assign n6154 = ~n5813 & ~n6153;
  assign n6155 = ~n5799 & n5813;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = pi02 & ~n6156;
  assign n6158 = ~pi02 & n6156;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = pi00 & ~n5813;
  assign n6161 = ~pi01 & n6160;
  assign n6162 = n6159 & ~n6161;
  assign n6163 = n6149 & n6162;
  assign n6164 = ~n5905 & ~n5921;
  assign n6165 = ~n5904 & ~n6164;
  assign n6166 = ~n5896 & ~n5926;
  assign n6167 = ~n6165 & n6166;
  assign n6168 = ~n5895 & ~n5947;
  assign n6169 = ~n6167 & n6168;
  assign n6170 = ~n5938 & ~n5946;
  assign n6171 = ~n6169 & n6170;
  assign n6172 = ~n5937 & ~n6171;
  assign n6173 = ~pi31 & ~n6172;
  assign n6174 = n5969 & ~n5979;
  assign n6175 = ~n5978 & ~n6174;
  assign n6176 = ~n5988 & n6175;
  assign n6177 = ~n5987 & ~n6176;
  assign n6178 = ~n5961 & n6177;
  assign n6179 = ~n5960 & ~n6178;
  assign n6180 = n5953 & n6179;
  assign n6181 = ~n6173 & ~n6180;
  assign n6182 = ~n6010 & n6021;
  assign n6183 = ~n6009 & ~n6019;
  assign n6184 = ~n6182 & n6183;
  assign n6185 = ~n6001 & ~n6018;
  assign n6186 = ~n6184 & n6185;
  assign n6187 = ~n6000 & ~n6186;
  assign n6188 = n5993 & n6187;
  assign n6189 = ~n6181 & ~n6188;
  assign n6190 = ~n6053 & n6061;
  assign n6191 = ~n6044 & ~n6052;
  assign n6192 = ~n6190 & n6191;
  assign n6193 = ~n6035 & ~n6043;
  assign n6194 = ~n6192 & n6193;
  assign n6195 = ~n6034 & ~n6194;
  assign n6196 = n6027 & n6195;
  assign n6197 = ~n6189 & ~n6196;
  assign n6198 = ~n6083 & n6092;
  assign n6199 = ~n6075 & ~n6084;
  assign n6200 = ~n6198 & n6199;
  assign n6201 = ~n6074 & ~n6102;
  assign n6202 = ~n6200 & n6201;
  assign n6203 = ~n6101 & ~n6202;
  assign n6204 = n6067 & n6203;
  assign n6205 = ~n6197 & ~n6204;
  assign n6206 = ~n6133 & ~n6141;
  assign n6207 = ~n6124 & ~n6132;
  assign n6208 = ~n6206 & n6207;
  assign n6209 = ~n6123 & ~n6208;
  assign n6210 = ~n6115 & ~n6209;
  assign n6211 = ~n6114 & ~n6210;
  assign n6212 = n6107 & n6211;
  assign n6213 = ~n6205 & ~n6212;
  assign n6214 = ~n5856 & n6157;
  assign n6215 = ~n5855 & ~n5864;
  assign n6216 = ~n6214 & n6215;
  assign n6217 = ~n5865 & ~n6216;
  assign n6218 = n6147 & n6217;
  assign n6219 = ~n6163 & ~n6218;
  assign n6220 = ~n6213 & n6219;
  assign n6221 = n84 & n6159;
  assign n6222 = n6149 & n6221;
  assign n6223 = ~n6220 & ~n6222;
  assign n6224 = ~n5848 & n6223;
  assign n6225 = ~n84 & ~n6161;
  assign n6226 = ~n6157 & ~n6225;
  assign n6227 = ~n6158 & ~n6226;
  assign n6228 = ~n5856 & n6227;
  assign n6229 = ~n5855 & ~n6228;
  assign n6230 = ~n5864 & n6229;
  assign n6231 = ~n5865 & ~n6230;
  assign n6232 = ~n6141 & ~n6231;
  assign n6233 = ~n6142 & ~n6232;
  assign n6234 = ~n6132 & n6233;
  assign n6235 = ~n6133 & ~n6234;
  assign n6236 = ~n6124 & ~n6235;
  assign n6237 = ~n6123 & ~n6236;
  assign n6238 = ~n6115 & ~n6237;
  assign n6239 = ~n6114 & ~n6238;
  assign n6240 = ~n6092 & ~n6239;
  assign n6241 = ~n6093 & ~n6240;
  assign n6242 = ~n6084 & ~n6241;
  assign n6243 = ~n6083 & ~n6242;
  assign n6244 = ~n6075 & ~n6243;
  assign n6245 = ~n6074 & ~n6244;
  assign n6246 = ~n6101 & ~n6245;
  assign n6247 = ~n6102 & ~n6246;
  assign n6248 = ~n6062 & ~n6247;
  assign n6249 = ~n6061 & ~n6248;
  assign n6250 = ~n6053 & ~n6249;
  assign n6251 = ~n6052 & ~n6250;
  assign n6252 = ~n6043 & ~n6251;
  assign n6253 = ~n6044 & ~n6252;
  assign n6254 = ~n6035 & ~n6253;
  assign n6255 = ~n6034 & ~n6254;
  assign n6256 = n6023 & ~n6255;
  assign n6257 = ~n6023 & n6255;
  assign n6258 = ~n6256 & ~n6257;
  assign n6259 = ~n6223 & n6258;
  assign n6260 = ~n6224 & ~n6259;
  assign n6261 = ~n5936 & n6223;
  assign n6262 = ~n6021 & ~n6255;
  assign n6263 = ~n6022 & ~n6262;
  assign n6264 = ~n6009 & ~n6263;
  assign n6265 = ~n6010 & ~n6264;
  assign n6266 = ~n6019 & ~n6265;
  assign n6267 = ~n6018 & ~n6266;
  assign n6268 = ~n6000 & ~n6267;
  assign n6269 = ~n6001 & ~n6268;
  assign n6270 = ~n5970 & ~n6269;
  assign n6271 = ~n5969 & ~n6270;
  assign n6272 = ~n5979 & ~n6271;
  assign n6273 = ~n5978 & ~n6272;
  assign n6274 = ~n5988 & n6273;
  assign n6275 = ~n5987 & ~n6274;
  assign n6276 = ~n5960 & ~n6275;
  assign n6277 = ~n5961 & ~n6276;
  assign n6278 = ~n5949 & ~n6277;
  assign n6279 = ~n5914 & ~n6278;
  assign n6280 = ~n5921 & ~n6279;
  assign n6281 = ~n5922 & ~n6280;
  assign n6282 = ~n5905 & ~n6281;
  assign n6283 = ~n5904 & ~n6282;
  assign n6284 = ~n5896 & ~n6283;
  assign n6285 = ~n5895 & ~n6284;
  assign n6286 = ~n5946 & ~n6285;
  assign n6287 = ~n5947 & ~n6286;
  assign n6288 = ~n5939 & ~n6287;
  assign n6289 = n5939 & n6287;
  assign n6290 = ~n6223 & ~n6288;
  assign n6291 = ~n6289 & n6290;
  assign n6292 = ~n6261 & ~n6291;
  assign n6293 = pi31 & ~n6292;
  assign n6294 = ~n5894 & n6223;
  assign n6295 = ~n5897 & ~n6283;
  assign n6296 = n5897 & n6283;
  assign n6297 = ~n6223 & ~n6295;
  assign n6298 = ~n6296 & n6297;
  assign n6299 = ~n6294 & ~n6298;
  assign n6300 = pi29 & ~n6299;
  assign n6301 = ~n5945 & n6223;
  assign n6302 = n5948 & ~n6285;
  assign n6303 = ~n5948 & n6285;
  assign n6304 = ~n6223 & ~n6302;
  assign n6305 = ~n6303 & n6304;
  assign n6306 = ~n6301 & ~n6305;
  assign n6307 = pi30 & n6306;
  assign n6308 = ~pi29 & n6299;
  assign n6309 = ~n5906 & ~n6281;
  assign n6310 = n5906 & n6281;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = ~n6223 & ~n6311;
  assign n6313 = ~n5903 & n6223;
  assign n6314 = ~n6312 & ~n6313;
  assign n6315 = ~pi28 & ~n6314;
  assign n6316 = pi28 & n6314;
  assign n6317 = ~n5920 & n6223;
  assign n6318 = ~n5923 & ~n6279;
  assign n6319 = n5923 & n6279;
  assign n6320 = ~n6223 & ~n6318;
  assign n6321 = ~n6319 & n6320;
  assign n6322 = ~n6317 & ~n6321;
  assign n6323 = pi27 & ~n6322;
  assign n6324 = n5913 & n6223;
  assign n6325 = ~n5914 & ~n5949;
  assign n6326 = ~n6277 & ~n6325;
  assign n6327 = n6277 & n6325;
  assign n6328 = ~n6223 & ~n6326;
  assign n6329 = ~n6327 & n6328;
  assign n6330 = ~n6324 & ~n6329;
  assign n6331 = ~pi26 & n6330;
  assign n6332 = ~pi27 & n6322;
  assign n6333 = pi26 & ~n6330;
  assign n6334 = ~n5959 & n6223;
  assign n6335 = n5962 & ~n6275;
  assign n6336 = ~n5962 & n6275;
  assign n6337 = ~n6223 & ~n6335;
  assign n6338 = ~n6336 & n6337;
  assign n6339 = ~n6334 & ~n6338;
  assign n6340 = pi25 & n6339;
  assign n6341 = ~pi25 & ~n6339;
  assign n6342 = ~n5986 & n6223;
  assign n6343 = n5989 & ~n6273;
  assign n6344 = ~n5989 & n6273;
  assign n6345 = ~n6223 & ~n6343;
  assign n6346 = ~n6344 & n6345;
  assign n6347 = ~n6342 & ~n6346;
  assign n6348 = ~pi24 & n6347;
  assign n6349 = ~n5977 & n6223;
  assign n6350 = n5980 & ~n6271;
  assign n6351 = ~n5980 & n6271;
  assign n6352 = ~n6223 & ~n6350;
  assign n6353 = ~n6351 & n6352;
  assign n6354 = ~n6349 & ~n6353;
  assign n6355 = pi23 & ~n6354;
  assign n6356 = pi24 & ~n6347;
  assign n6357 = ~n5968 & n6223;
  assign n6358 = n5971 & ~n6269;
  assign n6359 = ~n5971 & n6269;
  assign n6360 = ~n6223 & ~n6358;
  assign n6361 = ~n6359 & n6360;
  assign n6362 = ~n6357 & ~n6361;
  assign n6363 = ~pi22 & n6362;
  assign n6364 = ~pi23 & n6354;
  assign n6365 = pi22 & ~n6362;
  assign n6366 = ~n5999 & n6223;
  assign n6367 = n6002 & ~n6267;
  assign n6368 = ~n6002 & n6267;
  assign n6369 = ~n6223 & ~n6367;
  assign n6370 = ~n6368 & n6369;
  assign n6371 = ~n6366 & ~n6370;
  assign n6372 = pi21 & ~n6371;
  assign n6373 = ~n6017 & n6223;
  assign n6374 = n6020 & ~n6265;
  assign n6375 = ~n6020 & n6265;
  assign n6376 = ~n6223 & ~n6374;
  assign n6377 = ~n6375 & n6376;
  assign n6378 = ~n6373 & ~n6377;
  assign n6379 = ~pi20 & n6378;
  assign n6380 = ~pi21 & n6371;
  assign n6381 = pi20 & ~n6378;
  assign n6382 = ~n6008 & n6223;
  assign n6383 = n6011 & ~n6263;
  assign n6384 = ~n6011 & n6263;
  assign n6385 = ~n6223 & ~n6383;
  assign n6386 = ~n6384 & n6385;
  assign n6387 = ~n6382 & ~n6386;
  assign n6388 = pi19 & ~n6387;
  assign n6389 = ~pi18 & n6260;
  assign n6390 = ~pi19 & n6387;
  assign n6391 = pi18 & ~n6260;
  assign n6392 = n6033 & n6223;
  assign n6393 = n6036 & ~n6253;
  assign n6394 = ~n6036 & n6253;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n6223 & n6395;
  assign n6397 = ~n6392 & ~n6396;
  assign n6398 = pi17 & ~n6397;
  assign n6399 = ~n6042 & n6223;
  assign n6400 = n6045 & ~n6251;
  assign n6401 = ~n6045 & n6251;
  assign n6402 = ~n6400 & ~n6401;
  assign n6403 = ~n6223 & n6402;
  assign n6404 = ~n6399 & ~n6403;
  assign n6405 = ~pi16 & n6404;
  assign n6406 = ~pi17 & n6397;
  assign n6407 = ~n6051 & n6223;
  assign n6408 = n6054 & ~n6249;
  assign n6409 = ~n6054 & n6249;
  assign n6410 = ~n6408 & ~n6409;
  assign n6411 = ~n6223 & n6410;
  assign n6412 = ~n6407 & ~n6411;
  assign n6413 = pi15 & ~n6412;
  assign n6414 = ~pi15 & n6412;
  assign n6415 = ~n6060 & n6223;
  assign n6416 = n6063 & ~n6247;
  assign n6417 = ~n6063 & n6247;
  assign n6418 = ~n6416 & ~n6417;
  assign n6419 = ~n6223 & n6418;
  assign n6420 = ~n6415 & ~n6419;
  assign n6421 = pi14 & ~n6420;
  assign n6422 = ~n6100 & n6223;
  assign n6423 = n6103 & ~n6245;
  assign n6424 = ~n6103 & n6245;
  assign n6425 = ~n6423 & ~n6424;
  assign n6426 = ~n6223 & n6425;
  assign n6427 = ~n6422 & ~n6426;
  assign n6428 = ~pi13 & n6427;
  assign n6429 = ~pi14 & n6420;
  assign n6430 = pi13 & ~n6427;
  assign n6431 = ~n6073 & n6223;
  assign n6432 = n6076 & ~n6243;
  assign n6433 = ~n6076 & n6243;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = ~n6223 & n6434;
  assign n6436 = ~n6431 & ~n6435;
  assign n6437 = ~pi12 & n6436;
  assign n6438 = pi12 & ~n6436;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = ~n6082 & n6223;
  assign n6441 = n6085 & ~n6241;
  assign n6442 = ~n6085 & n6241;
  assign n6443 = ~n6441 & ~n6442;
  assign n6444 = ~n6223 & n6443;
  assign n6445 = ~n6440 & ~n6444;
  assign n6446 = pi11 & ~n6445;
  assign n6447 = ~pi11 & n6445;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n6131 & n6223;
  assign n6450 = ~n6134 & ~n6233;
  assign n6451 = n6134 & n6233;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = ~n6223 & n6452;
  assign n6454 = ~n6449 & ~n6453;
  assign n6455 = ~pi07 & n6454;
  assign n6456 = ~n6122 & n6223;
  assign n6457 = n6125 & ~n6235;
  assign n6458 = ~n6125 & n6235;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = ~n6223 & n6459;
  assign n6461 = ~n6456 & ~n6460;
  assign n6462 = ~pi08 & n6461;
  assign n6463 = pi07 & ~n6454;
  assign n6464 = ~n6143 & ~n6231;
  assign n6465 = n6143 & n6231;
  assign n6466 = ~n6464 & ~n6465;
  assign n6467 = ~n6223 & ~n6466;
  assign n6468 = n6140 & n6223;
  assign n6469 = ~n6467 & ~n6468;
  assign n6470 = pi06 & n6469;
  assign n6471 = ~pi06 & ~n6469;
  assign n6472 = ~n5863 & n6223;
  assign n6473 = n5866 & ~n6229;
  assign n6474 = ~n5866 & n6229;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~n6223 & n6475;
  assign n6477 = ~n6472 & ~n6476;
  assign n6478 = pi05 & ~n6477;
  assign n6479 = ~n6471 & n6478;
  assign n6480 = ~n6463 & ~n6470;
  assign n6481 = ~n6479 & n6480;
  assign n6482 = ~n6455 & ~n6462;
  assign n6483 = ~n6481 & n6482;
  assign n6484 = pi08 & ~n6461;
  assign n6485 = ~n6455 & ~n6463;
  assign n6486 = ~n6470 & ~n6471;
  assign n6487 = ~pi05 & n6477;
  assign n6488 = ~n6478 & ~n6487;
  assign n6489 = ~n6462 & ~n6484;
  assign n6490 = n6485 & n6486;
  assign n6491 = n6488 & n6489;
  assign n6492 = n6490 & n6491;
  assign n6493 = pi00 & ~n5807;
  assign n6494 = ~pi01 & ~n6493;
  assign n6495 = pi01 & n6493;
  assign n6496 = ~n6494 & ~n6495;
  assign n6497 = ~n6223 & ~n6496;
  assign n6498 = ~n6160 & n6223;
  assign n6499 = ~n6497 & ~n6498;
  assign n6500 = pi02 & ~n6499;
  assign n6501 = pi00 & ~n6223;
  assign n6502 = ~pi01 & n6501;
  assign n6503 = ~n6500 & n6502;
  assign n6504 = ~pi02 & n6499;
  assign n6505 = ~n5854 & n6223;
  assign n6506 = ~n5857 & ~n6227;
  assign n6507 = n5857 & n6227;
  assign n6508 = ~n6506 & ~n6507;
  assign n6509 = ~n6223 & n6508;
  assign n6510 = ~n6505 & ~n6509;
  assign n6511 = pi04 & ~n6510;
  assign n6512 = ~pi04 & n6510;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = ~n6156 & n6223;
  assign n6515 = ~n6159 & ~n6225;
  assign n6516 = n6159 & n6225;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = ~n6223 & n6517;
  assign n6519 = ~n6514 & ~n6518;
  assign n6520 = pi03 & ~n6519;
  assign n6521 = ~pi03 & n6519;
  assign n6522 = ~n6520 & ~n6521;
  assign n6523 = n6513 & n6522;
  assign n6524 = ~n6503 & ~n6504;
  assign n6525 = n6523 & n6524;
  assign n6526 = ~n6512 & n6520;
  assign n6527 = ~n6511 & ~n6526;
  assign n6528 = ~n6525 & n6527;
  assign n6529 = n6492 & ~n6528;
  assign n6530 = ~n6483 & ~n6484;
  assign n6531 = ~n6529 & n6530;
  assign n6532 = ~n6500 & ~n6504;
  assign n6533 = n84 & n6532;
  assign n6534 = n6523 & n6533;
  assign n6535 = n6492 & n6534;
  assign n6536 = ~n6531 & ~n6535;
  assign n6537 = ~n6113 & n6223;
  assign n6538 = n6116 & ~n6237;
  assign n6539 = ~n6116 & n6237;
  assign n6540 = ~n6538 & ~n6539;
  assign n6541 = ~n6223 & n6540;
  assign n6542 = ~n6537 & ~n6541;
  assign n6543 = ~pi09 & n6542;
  assign n6544 = pi09 & ~n6542;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = ~n6091 & n6223;
  assign n6547 = n6094 & ~n6239;
  assign n6548 = ~n6094 & n6239;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = ~n6223 & n6549;
  assign n6551 = ~n6546 & ~n6550;
  assign n6552 = pi10 & ~n6551;
  assign n6553 = ~pi10 & n6551;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = n6439 & n6448;
  assign n6556 = n6545 & n6554;
  assign n6557 = n6555 & n6556;
  assign n6558 = ~n6536 & n6557;
  assign n6559 = n6543 & ~n6552;
  assign n6560 = ~n6447 & ~n6553;
  assign n6561 = ~n6559 & n6560;
  assign n6562 = ~n6438 & ~n6446;
  assign n6563 = ~n6561 & n6562;
  assign n6564 = ~n6437 & ~n6563;
  assign n6565 = ~n6558 & n6564;
  assign n6566 = ~n6430 & ~n6565;
  assign n6567 = ~n6428 & ~n6429;
  assign n6568 = ~n6566 & n6567;
  assign n6569 = ~n6421 & ~n6568;
  assign n6570 = ~n6414 & ~n6569;
  assign n6571 = pi16 & ~n6404;
  assign n6572 = ~n6413 & ~n6571;
  assign n6573 = ~n6570 & n6572;
  assign n6574 = ~n6405 & ~n6406;
  assign n6575 = ~n6573 & n6574;
  assign n6576 = ~n6391 & ~n6398;
  assign n6577 = ~n6575 & n6576;
  assign n6578 = ~n6389 & ~n6390;
  assign n6579 = ~n6577 & n6578;
  assign n6580 = ~n6381 & ~n6388;
  assign n6581 = ~n6579 & n6580;
  assign n6582 = ~n6379 & ~n6380;
  assign n6583 = ~n6581 & n6582;
  assign n6584 = ~n6365 & ~n6372;
  assign n6585 = ~n6583 & n6584;
  assign n6586 = ~n6363 & ~n6364;
  assign n6587 = ~n6585 & n6586;
  assign n6588 = ~n6355 & ~n6356;
  assign n6589 = ~n6587 & n6588;
  assign n6590 = ~n6341 & ~n6348;
  assign n6591 = ~n6589 & n6590;
  assign n6592 = ~n6333 & ~n6340;
  assign n6593 = ~n6591 & n6592;
  assign n6594 = ~n6331 & ~n6332;
  assign n6595 = ~n6593 & n6594;
  assign n6596 = ~n6316 & ~n6323;
  assign n6597 = ~n6595 & n6596;
  assign n6598 = ~n6308 & ~n6315;
  assign n6599 = ~n6597 & n6598;
  assign n6600 = ~n6300 & ~n6307;
  assign n6601 = ~n6599 & n6600;
  assign n6602 = ~pi31 & n6292;
  assign n6603 = ~pi30 & ~n6306;
  assign n6604 = ~n6602 & ~n6603;
  assign n6605 = ~n6601 & n6604;
  assign n6606 = ~n6293 & ~n6605;
  assign n6607 = n6260 & ~n6606;
  assign n6608 = ~n6389 & ~n6391;
  assign n6609 = ~n84 & ~n6502;
  assign n6610 = ~n6504 & n6609;
  assign n6611 = ~n6500 & ~n6610;
  assign n6612 = ~n6521 & ~n6611;
  assign n6613 = ~n6520 & ~n6612;
  assign n6614 = ~n6512 & ~n6613;
  assign n6615 = ~n6511 & ~n6614;
  assign n6616 = ~n6487 & ~n6615;
  assign n6617 = ~n6478 & ~n6616;
  assign n6618 = ~n6471 & ~n6617;
  assign n6619 = ~n6470 & ~n6618;
  assign n6620 = ~n6455 & ~n6619;
  assign n6621 = ~n6463 & ~n6620;
  assign n6622 = ~n6462 & ~n6621;
  assign n6623 = ~n6484 & ~n6622;
  assign n6624 = ~n6543 & ~n6623;
  assign n6625 = ~n6544 & ~n6624;
  assign n6626 = ~n6553 & ~n6625;
  assign n6627 = ~n6552 & ~n6626;
  assign n6628 = ~n6447 & ~n6627;
  assign n6629 = ~n6446 & ~n6628;
  assign n6630 = ~n6437 & ~n6629;
  assign n6631 = ~n6438 & ~n6630;
  assign n6632 = ~n6428 & ~n6631;
  assign n6633 = ~n6430 & ~n6632;
  assign n6634 = ~n6429 & ~n6633;
  assign n6635 = ~n6421 & ~n6634;
  assign n6636 = ~n6414 & ~n6635;
  assign n6637 = ~n6413 & ~n6636;
  assign n6638 = ~n6571 & n6637;
  assign n6639 = ~n6405 & ~n6638;
  assign n6640 = ~n6406 & n6639;
  assign n6641 = ~n6398 & ~n6640;
  assign n6642 = ~n6608 & ~n6641;
  assign n6643 = n6608 & n6641;
  assign n6644 = n6606 & ~n6642;
  assign n6645 = ~n6643 & n6644;
  assign n6646 = ~n6607 & ~n6645;
  assign n6647 = pi19 & n6646;
  assign n6648 = ~n6397 & ~n6606;
  assign n6649 = ~n6398 & ~n6406;
  assign n6650 = ~n6639 & ~n6649;
  assign n6651 = n6639 & n6649;
  assign n6652 = n6606 & ~n6650;
  assign n6653 = ~n6651 & n6652;
  assign n6654 = ~n6648 & ~n6653;
  assign n6655 = ~pi18 & n6654;
  assign n6656 = ~pi19 & ~n6646;
  assign n6657 = ~n6647 & ~n6655;
  assign n6658 = ~n6656 & n6657;
  assign n6659 = ~n6647 & ~n6658;
  assign n6660 = n6306 & ~n6606;
  assign n6661 = ~n6307 & ~n6603;
  assign n6662 = ~n6389 & ~n6641;
  assign n6663 = ~n6391 & ~n6662;
  assign n6664 = ~n6390 & ~n6663;
  assign n6665 = ~n6388 & ~n6664;
  assign n6666 = ~n6379 & ~n6665;
  assign n6667 = ~n6381 & ~n6666;
  assign n6668 = ~n6380 & ~n6667;
  assign n6669 = ~n6372 & ~n6668;
  assign n6670 = ~n6363 & ~n6669;
  assign n6671 = ~n6365 & ~n6670;
  assign n6672 = ~n6364 & ~n6671;
  assign n6673 = ~n6355 & ~n6672;
  assign n6674 = ~n6348 & ~n6673;
  assign n6675 = ~n6356 & ~n6674;
  assign n6676 = ~n6341 & ~n6675;
  assign n6677 = ~n6340 & ~n6676;
  assign n6678 = ~n6331 & ~n6677;
  assign n6679 = ~n6333 & ~n6678;
  assign n6680 = ~n6332 & ~n6679;
  assign n6681 = ~n6323 & ~n6680;
  assign n6682 = ~n6315 & ~n6681;
  assign n6683 = ~n6316 & ~n6682;
  assign n6684 = ~n6308 & ~n6683;
  assign n6685 = ~n6300 & ~n6684;
  assign n6686 = n6661 & ~n6685;
  assign n6687 = ~n6661 & n6685;
  assign n6688 = n6606 & ~n6686;
  assign n6689 = ~n6687 & n6688;
  assign n6690 = ~n6660 & ~n6689;
  assign n6691 = ~pi31 & n6690;
  assign n6692 = n6292 & n6605;
  assign n6693 = ~n6307 & n6685;
  assign n6694 = ~n6603 & ~n6693;
  assign n6695 = ~n6602 & ~n6694;
  assign n6696 = n6602 & n6694;
  assign n6697 = n6606 & ~n6695;
  assign n6698 = ~n6696 & n6697;
  assign n6699 = ~n6691 & ~n6692;
  assign n6700 = ~n6698 & n6699;
  assign n6701 = pi31 & ~n6690;
  assign n6702 = ~n6299 & ~n6606;
  assign n6703 = ~n6300 & ~n6308;
  assign n6704 = n6683 & ~n6703;
  assign n6705 = ~n6683 & n6703;
  assign n6706 = n6606 & ~n6704;
  assign n6707 = ~n6705 & n6706;
  assign n6708 = ~n6702 & ~n6707;
  assign n6709 = pi30 & ~n6708;
  assign n6710 = ~n6701 & ~n6709;
  assign n6711 = ~n6314 & ~n6606;
  assign n6712 = ~n6315 & ~n6316;
  assign n6713 = ~n6681 & ~n6712;
  assign n6714 = n6681 & n6712;
  assign n6715 = n6606 & ~n6713;
  assign n6716 = ~n6714 & n6715;
  assign n6717 = ~n6711 & ~n6716;
  assign n6718 = pi29 & n6717;
  assign n6719 = n6322 & ~n6606;
  assign n6720 = ~n6323 & ~n6332;
  assign n6721 = ~n6679 & ~n6720;
  assign n6722 = n6679 & n6720;
  assign n6723 = n6606 & ~n6721;
  assign n6724 = ~n6722 & n6723;
  assign n6725 = ~n6719 & ~n6724;
  assign n6726 = pi28 & n6725;
  assign n6727 = ~n6718 & ~n6726;
  assign n6728 = ~n6339 & ~n6606;
  assign n6729 = ~n6340 & ~n6341;
  assign n6730 = ~n6675 & ~n6729;
  assign n6731 = n6675 & n6729;
  assign n6732 = n6606 & ~n6730;
  assign n6733 = ~n6731 & n6732;
  assign n6734 = ~n6728 & ~n6733;
  assign n6735 = ~pi26 & ~n6734;
  assign n6736 = ~pi30 & n6708;
  assign n6737 = ~pi29 & ~n6717;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = n6330 & ~n6606;
  assign n6740 = ~n6331 & ~n6333;
  assign n6741 = ~n6677 & ~n6740;
  assign n6742 = n6677 & n6740;
  assign n6743 = n6606 & ~n6741;
  assign n6744 = ~n6742 & n6743;
  assign n6745 = ~n6739 & ~n6744;
  assign n6746 = ~pi27 & ~n6745;
  assign n6747 = ~pi28 & ~n6725;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = pi27 & n6745;
  assign n6750 = pi26 & n6734;
  assign n6751 = ~n6735 & ~n6750;
  assign n6752 = ~n6749 & n6751;
  assign n6753 = n6748 & n6752;
  assign n6754 = n6727 & n6753;
  assign n6755 = n6738 & n6754;
  assign n6756 = n6710 & n6755;
  assign n6757 = n6700 & n6756;
  assign n6758 = n6347 & ~n6606;
  assign n6759 = ~n6348 & ~n6356;
  assign n6760 = ~n6673 & ~n6759;
  assign n6761 = n6673 & n6759;
  assign n6762 = n6606 & ~n6760;
  assign n6763 = ~n6761 & n6762;
  assign n6764 = ~n6758 & ~n6763;
  assign n6765 = pi25 & n6764;
  assign n6766 = ~pi25 & ~n6764;
  assign n6767 = n6354 & ~n6606;
  assign n6768 = ~n6355 & ~n6364;
  assign n6769 = ~n6671 & ~n6768;
  assign n6770 = n6671 & n6768;
  assign n6771 = n6606 & ~n6769;
  assign n6772 = ~n6770 & n6771;
  assign n6773 = ~n6767 & ~n6772;
  assign n6774 = pi24 & n6773;
  assign n6775 = ~pi24 & ~n6773;
  assign n6776 = n6362 & ~n6606;
  assign n6777 = ~n6363 & ~n6365;
  assign n6778 = ~n6669 & ~n6777;
  assign n6779 = n6669 & n6777;
  assign n6780 = n6606 & ~n6778;
  assign n6781 = ~n6779 & n6780;
  assign n6782 = ~n6776 & ~n6781;
  assign n6783 = ~pi23 & ~n6782;
  assign n6784 = pi23 & n6782;
  assign n6785 = n6371 & ~n6606;
  assign n6786 = ~n6372 & ~n6380;
  assign n6787 = ~n6667 & ~n6786;
  assign n6788 = n6667 & n6786;
  assign n6789 = n6606 & ~n6787;
  assign n6790 = ~n6788 & n6789;
  assign n6791 = ~n6785 & ~n6790;
  assign n6792 = pi22 & n6791;
  assign n6793 = ~n6784 & ~n6792;
  assign n6794 = ~pi22 & ~n6791;
  assign n6795 = ~n6783 & ~n6794;
  assign n6796 = n6793 & n6795;
  assign n6797 = ~n6774 & n6796;
  assign n6798 = ~n6775 & n6797;
  assign n6799 = ~n6765 & n6798;
  assign n6800 = ~n6766 & n6799;
  assign n6801 = n6757 & n6800;
  assign n6802 = ~n6378 & ~n6606;
  assign n6803 = ~n6379 & ~n6381;
  assign n6804 = n6665 & ~n6803;
  assign n6805 = ~n6665 & n6803;
  assign n6806 = n6606 & ~n6804;
  assign n6807 = ~n6805 & n6806;
  assign n6808 = ~n6802 & ~n6807;
  assign n6809 = ~pi21 & n6808;
  assign n6810 = pi21 & ~n6808;
  assign n6811 = ~n6387 & ~n6606;
  assign n6812 = ~n6388 & ~n6390;
  assign n6813 = n6663 & ~n6812;
  assign n6814 = ~n6663 & n6812;
  assign n6815 = n6606 & ~n6813;
  assign n6816 = ~n6814 & n6815;
  assign n6817 = ~n6811 & ~n6816;
  assign n6818 = pi20 & ~n6817;
  assign n6819 = ~n6810 & ~n6818;
  assign n6820 = ~pi20 & n6817;
  assign n6821 = ~n6809 & ~n6820;
  assign n6822 = n6819 & n6821;
  assign n6823 = n6801 & n6822;
  assign n6824 = ~n6659 & n6823;
  assign n6825 = ~n6809 & ~n6819;
  assign n6826 = n6801 & ~n6825;
  assign n6827 = ~n6783 & ~n6793;
  assign n6828 = ~n6774 & ~n6827;
  assign n6829 = ~n6775 & ~n6828;
  assign n6830 = ~n6766 & n6829;
  assign n6831 = ~n6765 & ~n6830;
  assign n6832 = n6757 & n6831;
  assign n6833 = n6735 & ~n6749;
  assign n6834 = n6748 & ~n6833;
  assign n6835 = n6727 & ~n6834;
  assign n6836 = n6738 & ~n6835;
  assign n6837 = n6710 & ~n6836;
  assign n6838 = n6700 & ~n6837;
  assign n6839 = ~n6832 & n6838;
  assign n6840 = ~n6801 & ~n6839;
  assign n6841 = ~n6826 & ~n6840;
  assign n6842 = ~n6824 & ~n6841;
  assign n6843 = pi18 & ~n6654;
  assign n6844 = n6658 & ~n6843;
  assign n6845 = n6823 & n6844;
  assign n6846 = ~n6404 & ~n6606;
  assign n6847 = ~n6405 & ~n6571;
  assign n6848 = n6637 & ~n6847;
  assign n6849 = ~n6637 & n6847;
  assign n6850 = ~n6848 & ~n6849;
  assign n6851 = n6606 & n6850;
  assign n6852 = ~n6846 & ~n6851;
  assign n6853 = pi17 & ~n6852;
  assign n6854 = ~n6413 & ~n6414;
  assign n6855 = ~n6635 & ~n6854;
  assign n6856 = n6635 & n6854;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = n6606 & ~n6857;
  assign n6859 = ~n6412 & ~n6606;
  assign n6860 = ~n6858 & ~n6859;
  assign n6861 = ~pi16 & n6860;
  assign n6862 = ~pi17 & n6852;
  assign n6863 = ~n6861 & ~n6862;
  assign n6864 = pi16 & ~n6860;
  assign n6865 = ~n6421 & ~n6429;
  assign n6866 = ~n6633 & ~n6865;
  assign n6867 = n6633 & n6865;
  assign n6868 = ~n6866 & ~n6867;
  assign n6869 = n6606 & ~n6868;
  assign n6870 = ~n6420 & ~n6606;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = ~pi15 & n6871;
  assign n6873 = ~n6864 & n6872;
  assign n6874 = ~n6428 & ~n6430;
  assign n6875 = ~n6631 & ~n6874;
  assign n6876 = n6631 & n6874;
  assign n6877 = ~n6875 & ~n6876;
  assign n6878 = n6606 & ~n6877;
  assign n6879 = ~n6427 & ~n6606;
  assign n6880 = ~n6878 & ~n6879;
  assign n6881 = pi14 & ~n6880;
  assign n6882 = pi15 & ~n6871;
  assign n6883 = ~n6864 & ~n6881;
  assign n6884 = ~n6882 & n6883;
  assign n6885 = n6863 & ~n6873;
  assign n6886 = ~n6884 & n6885;
  assign n6887 = ~n6853 & ~n6886;
  assign n6888 = n6845 & n6887;
  assign n6889 = ~n6842 & ~n6888;
  assign n6890 = ~n6445 & ~n6606;
  assign n6891 = n6448 & ~n6627;
  assign n6892 = ~n6448 & n6627;
  assign n6893 = ~n6891 & ~n6892;
  assign n6894 = n6606 & n6893;
  assign n6895 = ~n6890 & ~n6894;
  assign n6896 = ~pi12 & n6895;
  assign n6897 = ~n6551 & ~n6606;
  assign n6898 = n6554 & ~n6625;
  assign n6899 = ~n6554 & n6625;
  assign n6900 = ~n6898 & ~n6899;
  assign n6901 = n6606 & n6900;
  assign n6902 = ~n6897 & ~n6901;
  assign n6903 = pi11 & ~n6902;
  assign n6904 = n6469 & ~n6606;
  assign n6905 = n6486 & ~n6617;
  assign n6906 = ~n6486 & n6617;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = n6606 & n6907;
  assign n6909 = ~n6904 & ~n6908;
  assign n6910 = pi07 & ~n6909;
  assign n6911 = ~n6454 & ~n6606;
  assign n6912 = n6485 & ~n6619;
  assign n6913 = ~n6485 & n6619;
  assign n6914 = ~n6912 & ~n6913;
  assign n6915 = n6606 & n6914;
  assign n6916 = ~n6911 & ~n6915;
  assign n6917 = pi08 & ~n6916;
  assign n6918 = ~pi07 & n6909;
  assign n6919 = ~n6477 & ~n6606;
  assign n6920 = n6488 & ~n6615;
  assign n6921 = ~n6488 & n6615;
  assign n6922 = ~n6920 & ~n6921;
  assign n6923 = n6606 & n6922;
  assign n6924 = ~n6919 & ~n6923;
  assign n6925 = ~pi06 & n6924;
  assign n6926 = pi06 & ~n6924;
  assign n6927 = ~n6510 & ~n6606;
  assign n6928 = n6513 & ~n6613;
  assign n6929 = ~n6513 & n6613;
  assign n6930 = ~n6928 & ~n6929;
  assign n6931 = n6606 & n6930;
  assign n6932 = ~n6927 & ~n6931;
  assign n6933 = pi05 & ~n6932;
  assign n6934 = ~pi05 & n6932;
  assign n6935 = ~n6519 & ~n6606;
  assign n6936 = n6522 & ~n6611;
  assign n6937 = ~n6522 & n6611;
  assign n6938 = ~n6936 & ~n6937;
  assign n6939 = n6606 & n6938;
  assign n6940 = ~n6935 & ~n6939;
  assign n6941 = ~pi04 & n6940;
  assign n6942 = ~n6532 & n6609;
  assign n6943 = n6532 & ~n6609;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = n6606 & ~n6944;
  assign n6946 = ~n6499 & ~n6606;
  assign n6947 = ~n6945 & ~n6946;
  assign n6948 = pi03 & ~n6947;
  assign n6949 = pi04 & ~n6940;
  assign n6950 = pi00 & ~n6220;
  assign n6951 = ~pi01 & ~n6950;
  assign n6952 = pi01 & n6950;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = n6606 & n6953;
  assign n6955 = n6501 & ~n6606;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = pi02 & n6956;
  assign n6958 = pi00 & ~n6606;
  assign n6959 = ~pi01 & ~n6958;
  assign n6960 = ~n6957 & n6959;
  assign n6961 = ~pi03 & n6947;
  assign n6962 = ~pi02 & ~n6956;
  assign n6963 = ~n6961 & ~n6962;
  assign n6964 = ~n6960 & n6963;
  assign n6965 = ~n6948 & ~n6949;
  assign n6966 = ~n6964 & n6965;
  assign n6967 = ~n6934 & ~n6941;
  assign n6968 = ~n6966 & n6967;
  assign n6969 = ~n6926 & ~n6933;
  assign n6970 = ~n6968 & n6969;
  assign n6971 = ~n6918 & ~n6925;
  assign n6972 = ~n6970 & n6971;
  assign n6973 = ~n6910 & ~n6917;
  assign n6974 = ~n6972 & n6973;
  assign n6975 = ~n6461 & ~n6606;
  assign n6976 = n6489 & ~n6621;
  assign n6977 = ~n6489 & n6621;
  assign n6978 = ~n6976 & ~n6977;
  assign n6979 = n6606 & n6978;
  assign n6980 = ~n6975 & ~n6979;
  assign n6981 = ~pi09 & n6980;
  assign n6982 = ~pi08 & n6916;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = ~n6974 & n6983;
  assign n6985 = ~n6542 & ~n6606;
  assign n6986 = n6545 & ~n6623;
  assign n6987 = ~n6545 & n6623;
  assign n6988 = ~n6986 & ~n6987;
  assign n6989 = n6606 & n6988;
  assign n6990 = ~n6985 & ~n6989;
  assign n6991 = pi10 & ~n6990;
  assign n6992 = ~n6439 & ~n6629;
  assign n6993 = n6439 & n6629;
  assign n6994 = ~n6992 & ~n6993;
  assign n6995 = n6606 & ~n6994;
  assign n6996 = ~n6436 & ~n6606;
  assign n6997 = ~n6995 & ~n6996;
  assign n6998 = ~pi13 & n6997;
  assign n6999 = pi09 & ~n6980;
  assign n7000 = ~n6991 & ~n6998;
  assign n7001 = ~n6999 & n7000;
  assign n7002 = ~n6984 & n7001;
  assign n7003 = ~pi11 & n6902;
  assign n7004 = ~pi10 & n6990;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = ~n7002 & n7005;
  assign n7007 = ~n6903 & ~n7006;
  assign n7008 = ~n6896 & ~n7007;
  assign n7009 = pi13 & ~n6997;
  assign n7010 = pi12 & ~n6895;
  assign n7011 = ~n7009 & ~n7010;
  assign n7012 = ~n7008 & n7011;
  assign n7013 = ~pi14 & n6880;
  assign n7014 = ~n6853 & ~n6872;
  assign n7015 = ~n6998 & ~n7013;
  assign n7016 = n7014 & n7015;
  assign n7017 = n6863 & n7016;
  assign n7018 = n6884 & n7017;
  assign n7019 = ~n7012 & n7018;
  assign n7020 = n6845 & n7019;
  assign n7021 = ~pi06 & ~pi13;
  assign n7022 = ~pi14 & ~pi21;
  assign n7023 = n7021 & n7022;
  assign n7024 = n65 & n91;
  assign n7025 = n94 & n7024;
  assign n7026 = n79 & n7023;
  assign n7027 = n89 & n7026;
  assign n7028 = n86 & n7025;
  assign n7029 = n7027 & n7028;
  assign n7030 = n74 & n7029;
  assign n7031 = ~n7020 & ~n7030;
  assign po00 = ~n6889 & n7031;
  assign po01 = n6606 & ~n7030;
  assign po02 = ~n6223 & ~n7030;
  assign po03 = ~n5813 & ~n7030;
  assign po04 = ~n5419 & ~n7030;
  assign po05 = ~n5037 & ~n7030;
  assign po06 = ~n4669 & ~n7030;
  assign po07 = ~n4317 & ~n7030;
  assign po08 = ~n3973 & ~n7030;
  assign po09 = ~n3646 & ~n7030;
  assign po10 = ~n3338 & ~n7030;
  assign po11 = ~n3038 & ~n7030;
  assign po12 = ~n2756 & ~n7030;
  assign po13 = ~n2488 & ~n7030;
  assign po14 = ~n2230 & ~n7030;
  assign po15 = ~n1988 & ~n7030;
  assign po16 = ~n1761 & ~n7030;
  assign po17 = ~n1545 & ~n7030;
  assign po18 = ~n1347 & ~n7030;
  assign po19 = ~n1161 & ~n7030;
  assign po20 = ~n987 & ~n7030;
  assign po21 = ~n831 & ~n7030;
  assign po22 = ~n691 & ~n7030;
  assign po23 = ~n560 & ~n7030;
  assign po24 = ~n443 & ~n7030;
  assign po25 = ~n340 & ~n7030;
  assign po26 = ~n254 & ~n7030;
  assign po27 = ~n182 & ~n7030;
  assign po28 = ~n126 & ~n7030;
  assign po29 = n115 & ~n7030;
  assign n7062 = ~n84 & ~n109;
  assign n7063 = n101 & ~n7030;
  assign po30 = ~n7062 & n7063;
  assign n7065 = ~pi00 & ~pi02;
  assign po31 = n7063 & n7065;
endmodule


