// Benchmark "table_out_0_93" written by ABC on Wed Apr 26 17:06:20 2017

module table_out_0_93 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83,
    po84, po85, po86, po87, po88, po89, po90, po91, po92, po93  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82,
    po83, po84, po85, po86, po87, po88, po89, po90, po91, po92, po93;
  wire n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n238, n239, n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
    n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3487, n3488, n3489, n3490, n3491,
    n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
    n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
    n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
    n3593, n3594, n3595, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3725, n3726, n3727, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
    n3756, n3757, n3758, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4241, n4242,
    n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
    n4273, n4274, n4275, n4278, n4279, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4319, n4320, n4321, n4322, n4323, n4324, n4326, n4327,
    n4328, n4330, n4331, n4333, n4334, n4335, n4337, n4338, n4339, n4340,
    n4342, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
    n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
    n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
    n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
    n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
    n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
    n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
    n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
    n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4743, n4744,
    n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4823, n4824, n4825,
    n4826, n4827, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
    n4839, n4840, n4841, n4843, n4844, n4846, n4847, n4849, n4850, n4851,
    n4853, n4854, n4856, n4858, n4859, n4860, n4861, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
    n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
    n4907, n4908, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4955, n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
    n5016, n5017, n5018, n5019, n5022, n5023, n5024, n5025, n5026, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
    n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
    n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
    n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
    n5292, n5293, n5294, n5295, n5297, n5298, n5299, n5301, n5302, n5303,
    n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
    n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5472, n5473, n5474, n5475, n5476, n5477, n5479,
    n5480, n5481, n5484, n5485, n5486, n5487, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5543, n5544, n5547;
  assign n223 = pi044 & pi045;
  assign n224 = pi122 & ~n223;
  assign n225 = pi002 & ~pi003;
  assign n226 = pi000 & ~pi127;
  assign n227 = n225 & n226;
  assign n228 = ~pi001 & n227;
  assign n229 = ~pi004 & pi005;
  assign n230 = pi006 & n229;
  assign n231 = ~pi007 & n230;
  assign n232 = n228 & n231;
  assign n233 = ~pi012 & ~pi013;
  assign n234 = pi014 & ~pi015;
  assign n235 = n233 & n234;
  assign n236 = n232 & n235;
  assign po00 = n224 & n236;
  assign n238 = ~pi002 & pi003;
  assign n239 = n226 & n238;
  assign n240 = pi001 & n239;
  assign n241 = pi007 & n230;
  assign n242 = ~pi115 & n241;
  assign n243 = n240 & n242;
  assign n244 = ~pi007 & n240;
  assign n245 = n229 & n244;
  assign n246 = ~n243 & ~n245;
  assign n247 = ~pi112 & ~n246;
  assign n248 = pi035 & ~pi123;
  assign n249 = n247 & ~n248;
  assign n250 = ~pi005 & pi006;
  assign n251 = ~pi004 & n250;
  assign n252 = ~pi112 & n251;
  assign n253 = ~pi046 & n252;
  assign n254 = n244 & n253;
  assign n255 = ~pi079 & n254;
  assign n256 = ~pi031 & n255;
  assign n257 = ~n249 & ~n256;
  assign n258 = ~pi056 & pi122;
  assign n259 = pi055 & n258;
  assign n260 = ~pi044 & pi055;
  assign n261 = n224 & ~n260;
  assign n262 = ~n259 & ~n261;
  assign n263 = pi123 & ~n247;
  assign n264 = ~n262 & ~n263;
  assign n265 = pi122 & ~n264;
  assign n266 = ~n257 & ~n265;
  assign n267 = ~pi019 & ~pi022;
  assign n268 = pi004 & pi005;
  assign n269 = ~pi006 & n268;
  assign n270 = ~pi018 & ~pi021;
  assign n271 = n269 & n270;
  assign n272 = n267 & n271;
  assign n273 = ~pi017 & pi020;
  assign n274 = pi001 & pi007;
  assign n275 = n227 & n274;
  assign n276 = pi016 & n275;
  assign n277 = n273 & n276;
  assign n278 = ~pi023 & n277;
  assign n279 = pi122 & n278;
  assign n280 = n272 & n279;
  assign n281 = ~n223 & n280;
  assign n282 = ~pi024 & ~pi025;
  assign n283 = ~pi027 & n282;
  assign n284 = ~pi026 & n283;
  assign n285 = pi112 & n284;
  assign n286 = ~pi123 & n285;
  assign n287 = n243 & n286;
  assign n288 = pi112 & n251;
  assign n289 = pi002 & pi003;
  assign n290 = n226 & n289;
  assign n291 = pi001 & n290;
  assign n292 = ~pi007 & n291;
  assign n293 = pi061 & n292;
  assign n294 = n288 & n293;
  assign n295 = ~pi035 & ~pi123;
  assign n296 = pi112 & n244;
  assign n297 = n295 & n296;
  assign n298 = n229 & n297;
  assign n299 = ~n294 & ~n298;
  assign n300 = ~n287 & n299;
  assign n301 = ~n281 & n300;
  assign n302 = pi122 & n262;
  assign n303 = pi123 & n255;
  assign n304 = pi001 & ~pi007;
  assign n305 = n227 & n304;
  assign n306 = n250 & n305;
  assign n307 = n244 & n269;
  assign n308 = ~pi005 & pi007;
  assign n309 = ~pi004 & n308;
  assign n310 = n240 & n309;
  assign n311 = ~n307 & ~n310;
  assign n312 = ~n306 & n311;
  assign n313 = ~n303 & n312;
  assign n314 = ~n302 & ~n313;
  assign n315 = pi007 & n291;
  assign n316 = ~pi004 & ~pi005;
  assign n317 = ~pi006 & n316;
  assign n318 = n315 & n317;
  assign n319 = ~pi061 & ~pi065;
  assign n320 = n252 & n291;
  assign n321 = ~n319 & n320;
  assign n322 = ~n318 & ~n321;
  assign n323 = ~n302 & ~n322;
  assign n324 = ~pi122 & n288;
  assign n325 = n315 & n324;
  assign n326 = ~n323 & ~n325;
  assign n327 = ~n314 & n326;
  assign n328 = n301 & n327;
  assign po01 = n266 | ~n328;
  assign n330 = pi079 & n254;
  assign n331 = ~n302 & n330;
  assign n332 = ~pi009 & ~pi010;
  assign n333 = pi012 & pi013;
  assign n334 = ~pi011 & n333;
  assign n335 = n332 & n334;
  assign n336 = pi005 & ~pi006;
  assign n337 = ~pi004 & n336;
  assign n338 = n275 & n337;
  assign n339 = ~pi008 & pi014;
  assign n340 = n338 & n339;
  assign n341 = n335 & n340;
  assign n342 = pi004 & pi006;
  assign n343 = ~pi005 & n342;
  assign n344 = n240 & n343;
  assign n345 = pi004 & ~pi005;
  assign n346 = ~pi006 & n345;
  assign n347 = n239 & n274;
  assign n348 = ~pi112 & n347;
  assign n349 = n346 & n348;
  assign n350 = ~n344 & ~n349;
  assign n351 = ~n341 & n350;
  assign n352 = ~pi025 & ~pi026;
  assign n353 = ~pi024 & n352;
  assign n354 = pi027 & n353;
  assign n355 = ~n351 & n354;
  assign n356 = ~n302 & n355;
  assign n357 = pi011 & ~pi012;
  assign n358 = ~pi013 & n357;
  assign n359 = n332 & n358;
  assign n360 = n284 & n359;
  assign n361 = ~pi008 & n234;
  assign n362 = n338 & n361;
  assign n363 = ~pi047 & n362;
  assign n364 = n360 & n363;
  assign n365 = ~n262 & n364;
  assign n366 = ~n356 & ~n365;
  assign po02 = n331 | ~n366;
  assign n368 = pi017 & pi020;
  assign n369 = n276 & n368;
  assign n370 = ~pi023 & n369;
  assign n371 = n272 & n370;
  assign n372 = n273 & n275;
  assign n373 = ~pi016 & n372;
  assign n374 = pi018 & pi021;
  assign n375 = pi019 & pi022;
  assign n376 = n374 & n375;
  assign n377 = ~pi023 & n376;
  assign n378 = n373 & n377;
  assign n379 = n230 & n378;
  assign n380 = ~n371 & ~n379;
  assign n381 = ~n284 & ~n380;
  assign n382 = pi044 & pi122;
  assign n383 = pi045 & n382;
  assign n384 = ~pi023 & n230;
  assign n385 = ~pi019 & pi022;
  assign n386 = n384 & n385;
  assign n387 = ~pi018 & pi021;
  assign n388 = n373 & n387;
  assign n389 = n386 & n388;
  assign n390 = ~n383 & n389;
  assign n391 = ~pi016 & n275;
  assign n392 = ~pi017 & n391;
  assign n393 = n376 & n392;
  assign n394 = pi023 & n230;
  assign n395 = n393 & n394;
  assign n396 = pi020 & n395;
  assign n397 = ~n223 & n396;
  assign n398 = ~n390 & ~n397;
  assign n399 = ~pi005 & ~pi006;
  assign n400 = n275 & n399;
  assign n401 = ~n302 & n400;
  assign n402 = n398 & ~n401;
  assign n403 = ~n381 & n402;
  assign n404 = ~pi026 & ~pi027;
  assign n405 = ~pi023 & n343;
  assign n406 = ~n404 & n405;
  assign n407 = ~pi020 & n391;
  assign n408 = ~pi017 & n407;
  assign n409 = ~pi022 & n374;
  assign n410 = n408 & n409;
  assign n411 = ~pi019 & n410;
  assign n412 = n406 & n411;
  assign n413 = ~po00 & ~n412;
  assign n414 = ~pi001 & ~pi007;
  assign n415 = n251 & n414;
  assign n416 = n290 & n415;
  assign n417 = pi008 & n416;
  assign n418 = n332 & n417;
  assign n419 = n358 & n418;
  assign n420 = ~n404 & n419;
  assign n421 = ~pi014 & n420;
  assign n422 = pi015 & n421;
  assign n423 = n345 & ~n383;
  assign n424 = ~pi006 & pi007;
  assign n425 = n291 & n354;
  assign n426 = ~n424 & n425;
  assign n427 = n423 & n426;
  assign n428 = pi061 & n427;
  assign n429 = ~n422 & ~n428;
  assign n430 = n413 & n429;
  assign po03 = ~n403 | ~n430;
  assign n432 = n251 & ~n383;
  assign n433 = pi022 & pi023;
  assign n434 = pi017 & ~pi020;
  assign n435 = n276 & n434;
  assign n436 = ~pi019 & n435;
  assign n437 = ~pi018 & n436;
  assign n438 = n433 & n437;
  assign n439 = ~pi001 & n239;
  assign n440 = ~n411 & ~n439;
  assign n441 = ~n438 & n440;
  assign n442 = n432 & ~n441;
  assign n443 = ~n383 & n405;
  assign n444 = n435 & n443;
  assign n445 = n374 & n444;
  assign n446 = pi021 & n433;
  assign n447 = pi018 & n435;
  assign n448 = n343 & n447;
  assign n449 = n446 & n448;
  assign n450 = pi020 & n405;
  assign n451 = pi018 & ~pi021;
  assign n452 = pi017 & n276;
  assign n453 = n451 & n452;
  assign n454 = n450 & n453;
  assign n455 = ~n449 & ~n454;
  assign n456 = ~n383 & ~n455;
  assign n457 = ~n445 & ~n456;
  assign n458 = pi014 & pi015;
  assign n459 = ~pi002 & ~pi003;
  assign n460 = n226 & n459;
  assign n461 = n304 & n460;
  assign n462 = pi012 & ~pi013;
  assign n463 = n461 & n462;
  assign n464 = n458 & n463;
  assign n465 = n337 & n464;
  assign n466 = n457 & ~n465;
  assign n467 = pi018 & pi022;
  assign n468 = n275 & n368;
  assign n469 = ~pi016 & n468;
  assign n470 = n467 & n469;
  assign n471 = n391 & n434;
  assign n472 = pi019 & ~pi022;
  assign n473 = n387 & n472;
  assign n474 = n471 & n473;
  assign n475 = ~n470 & ~n474;
  assign n476 = ~pi018 & n375;
  assign n477 = n471 & n476;
  assign n478 = n475 & ~n477;
  assign n479 = n443 & ~n478;
  assign n480 = n269 & ~n383;
  assign n481 = n228 & n480;
  assign n482 = n375 & n387;
  assign n483 = n343 & ~n383;
  assign n484 = pi023 & n471;
  assign n485 = n483 & n484;
  assign n486 = n482 & n485;
  assign n487 = ~n481 & ~n486;
  assign n488 = ~n479 & n487;
  assign n489 = n466 & n488;
  assign n490 = n373 & ~n383;
  assign n491 = n270 & n385;
  assign n492 = n230 & n491;
  assign n493 = n490 & n492;
  assign n494 = ~pi000 & ~pi127;
  assign n495 = n459 & n494;
  assign n496 = n304 & n495;
  assign n497 = n316 & n496;
  assign n498 = ~n383 & n497;
  assign n499 = ~n493 & ~n498;
  assign n500 = n436 & n451;
  assign n501 = n483 & n500;
  assign n502 = pi022 & n451;
  assign n503 = n483 & n502;
  assign n504 = n435 & n503;
  assign n505 = ~n501 & ~n504;
  assign n506 = pi023 & ~n505;
  assign n507 = n499 & ~n506;
  assign n508 = ~pi008 & ~pi014;
  assign n509 = n416 & n508;
  assign n510 = pi009 & pi010;
  assign n511 = pi011 & pi012;
  assign n512 = ~pi015 & n511;
  assign n513 = n510 & n512;
  assign n514 = n509 & n513;
  assign n515 = ~pi014 & pi015;
  assign n516 = ~pi008 & n515;
  assign n517 = n416 & n516;
  assign n518 = ~pi012 & pi013;
  assign n519 = ~pi011 & n518;
  assign n520 = n332 & n519;
  assign n521 = n517 & n520;
  assign n522 = ~n514 & ~n521;
  assign n523 = pi101 & pi103;
  assign n524 = ~pi102 & n523;
  assign n525 = ~n352 & n383;
  assign n526 = n524 & ~n525;
  assign n527 = ~n522 & ~n526;
  assign n528 = ~pi045 & n230;
  assign n529 = pi115 & n347;
  assign n530 = ~pi056 & n284;
  assign n531 = n529 & n530;
  assign n532 = n528 & n531;
  assign n533 = n230 & n284;
  assign n534 = ~pi044 & pi045;
  assign n535 = pi056 & n534;
  assign n536 = n533 & n535;
  assign n537 = n529 & n536;
  assign n538 = ~n532 & ~n537;
  assign n539 = ~n527 & n538;
  assign n540 = pi023 & n251;
  assign n541 = pi020 & n540;
  assign n542 = n392 & n541;
  assign n543 = pi022 & n374;
  assign n544 = n542 & n543;
  assign n545 = ~n383 & n544;
  assign n546 = n337 & n461;
  assign n547 = pi013 & pi015;
  assign n548 = pi014 & n547;
  assign n549 = n546 & n548;
  assign n550 = ~n545 & ~n549;
  assign n551 = ~pi023 & n432;
  assign n552 = ~pi018 & pi022;
  assign n553 = pi019 & ~pi021;
  assign n554 = ~n552 & n553;
  assign n555 = n471 & n554;
  assign n556 = n551 & n555;
  assign n557 = n374 & n385;
  assign n558 = n471 & n557;
  assign n559 = n480 & n558;
  assign n560 = n304 & n494;
  assign n561 = ~n383 & n560;
  assign n562 = ~n459 & n561;
  assign n563 = n317 & n562;
  assign n564 = ~n559 & ~n563;
  assign n565 = ~n556 & n564;
  assign n566 = n550 & n565;
  assign n567 = n539 & n566;
  assign n568 = n507 & n567;
  assign n569 = n267 & n374;
  assign n570 = n343 & n373;
  assign n571 = n569 & n570;
  assign n572 = ~n383 & n571;
  assign n573 = n290 & n414;
  assign n574 = pi005 & n342;
  assign n575 = n573 & n574;
  assign n576 = ~n383 & n575;
  assign n577 = ~n572 & ~n576;
  assign n578 = ~pi039 & ~n577;
  assign n579 = pi009 & ~pi010;
  assign n580 = n338 & n508;
  assign n581 = n579 & n580;
  assign n582 = ~pi015 & n581;
  assign n583 = ~n383 & n582;
  assign n584 = ~pi011 & ~n233;
  assign n585 = n583 & n584;
  assign n586 = pi023 & ~n383;
  assign n587 = pi020 & n251;
  assign n588 = n586 & n587;
  assign n589 = n452 & n588;
  assign n590 = n491 & n589;
  assign n591 = ~pi004 & pi006;
  assign n592 = ~pi001 & pi007;
  assign n593 = n239 & n592;
  assign n594 = n591 & n593;
  assign n595 = ~n383 & n594;
  assign n596 = pi005 & n595;
  assign n597 = n229 & ~n383;
  assign n598 = n439 & n597;
  assign n599 = ~pi007 & n598;
  assign n600 = ~n596 & ~n599;
  assign n601 = ~n590 & n600;
  assign n602 = ~n585 & n601;
  assign n603 = ~n578 & n602;
  assign n604 = n568 & n603;
  assign n605 = n489 & n604;
  assign n606 = ~n442 & n605;
  assign n607 = n354 & n496;
  assign n608 = n574 & n607;
  assign n609 = ~pi023 & n251;
  assign n610 = n557 & n609;
  assign n611 = n354 & n408;
  assign n612 = n610 & n611;
  assign n613 = ~n608 & ~n612;
  assign n614 = ~n383 & ~n613;
  assign n615 = pi031 & n255;
  assign n616 = n295 & n615;
  assign n617 = n354 & n616;
  assign n618 = pi026 & n282;
  assign n619 = ~pi027 & n618;
  assign n620 = ~pi013 & n514;
  assign n621 = n619 & n620;
  assign n622 = n524 & n621;
  assign n623 = ~n617 & ~n622;
  assign n624 = ~n614 & n623;
  assign n625 = n290 & n592;
  assign n626 = n408 & n451;
  assign n627 = n472 & n626;
  assign n628 = pi023 & n627;
  assign n629 = ~n625 & ~n628;
  assign n630 = n343 & ~n629;
  assign n631 = n354 & n630;
  assign n632 = n373 & n609;
  assign n633 = n557 & n632;
  assign n634 = n619 & n633;
  assign n635 = n378 & n432;
  assign n636 = ~n634 & ~n635;
  assign n637 = n292 & n399;
  assign n638 = ~pi004 & n637;
  assign n639 = n619 & n638;
  assign n640 = n636 & ~n639;
  assign n641 = ~n631 & n640;
  assign n642 = n624 & n641;
  assign n643 = n392 & n557;
  assign n644 = ~pi020 & n643;
  assign n645 = n405 & n644;
  assign n646 = ~n404 & n645;
  assign n647 = n224 & n232;
  assign n648 = pi014 & n233;
  assign n649 = n647 & n648;
  assign n650 = pi015 & n649;
  assign n651 = n377 & n570;
  assign n652 = n619 & n651;
  assign n653 = ~n650 & ~n652;
  assign n654 = ~pi014 & ~pi015;
  assign n655 = n420 & n654;
  assign n656 = n653 & ~n655;
  assign n657 = ~n646 & n656;
  assign n658 = ~pi061 & n427;
  assign n659 = n239 & n414;
  assign n660 = n317 & n659;
  assign n661 = ~pi017 & n276;
  assign n662 = n270 & n661;
  assign n663 = n472 & n662;
  assign n664 = ~pi020 & n663;
  assign n665 = n405 & n664;
  assign n666 = ~n660 & ~n665;
  assign n667 = ~n404 & ~n666;
  assign n668 = ~n658 & ~n667;
  assign n669 = n657 & n668;
  assign n670 = n642 & n669;
  assign po04 = ~n606 | ~n670;
  assign n672 = n387 & n392;
  assign n673 = ~n375 & n672;
  assign n674 = n480 & n673;
  assign n675 = n269 & n305;
  assign n676 = pi016 & n675;
  assign n677 = n434 & n676;
  assign n678 = n267 & n387;
  assign n679 = n677 & n678;
  assign n680 = pi072 & n679;
  assign n681 = n505 & ~n680;
  assign n682 = ~n674 & n681;
  assign n683 = ~pi031 & ~pi034;
  assign n684 = ~pi012 & n654;
  assign n685 = n317 & n460;
  assign n686 = n304 & n685;
  assign n687 = pi013 & n686;
  assign n688 = n684 & n687;
  assign n689 = n227 & n592;
  assign n690 = n230 & n689;
  assign n691 = n518 & n690;
  assign n692 = n654 & n691;
  assign n693 = ~n688 & ~n692;
  assign n694 = n241 & n495;
  assign n695 = pi001 & n694;
  assign n696 = pi039 & n695;
  assign n697 = n693 & ~n696;
  assign n698 = n683 & ~n697;
  assign n699 = n251 & n625;
  assign n700 = n579 & n699;
  assign n701 = pi008 & n700;
  assign n702 = ~pi013 & n511;
  assign n703 = n701 & n702;
  assign n704 = pi008 & ~pi014;
  assign n705 = pi011 & pi013;
  assign n706 = ~pi001 & n290;
  assign n707 = n251 & n706;
  assign n708 = pi007 & pi009;
  assign n709 = pi010 & n708;
  assign n710 = n707 & n709;
  assign n711 = n705 & n710;
  assign n712 = n704 & n711;
  assign n713 = pi015 & n712;
  assign n714 = ~n703 & ~n713;
  assign n715 = ~n698 & n714;
  assign n716 = ~n283 & ~n353;
  assign n717 = ~n404 & ~n716;
  assign n718 = n651 & n717;
  assign n719 = ~pi023 & n679;
  assign n720 = ~n718 & ~n719;
  assign n721 = n715 & n720;
  assign n722 = n682 & n721;
  assign n723 = n394 & n409;
  assign n724 = n436 & n723;
  assign n725 = n369 & n384;
  assign n726 = n385 & n387;
  assign n727 = n725 & n726;
  assign n728 = ~n724 & ~n727;
  assign n729 = pi021 & n385;
  assign n730 = n275 & n434;
  assign n731 = n394 & n730;
  assign n732 = pi016 & n731;
  assign n733 = n729 & n732;
  assign n734 = n230 & n452;
  assign n735 = ~pi020 & n734;
  assign n736 = ~pi018 & ~pi019;
  assign n737 = ~pi022 & n736;
  assign n738 = ~pi021 & n385;
  assign n739 = ~n737 & ~n738;
  assign n740 = n735 & ~n739;
  assign n741 = n230 & n277;
  assign n742 = n726 & n741;
  assign n743 = ~n740 & ~n742;
  assign n744 = ~n733 & n743;
  assign n745 = n728 & n744;
  assign n746 = pi017 & n675;
  assign n747 = ~pi016 & n746;
  assign n748 = ~pi018 & n385;
  assign n749 = ~pi020 & ~pi023;
  assign n750 = n748 & n749;
  assign n751 = n747 & n750;
  assign n752 = pi021 & n736;
  assign n753 = pi022 & ~pi023;
  assign n754 = n752 & n753;
  assign n755 = pi020 & n747;
  assign n756 = n754 & n755;
  assign n757 = ~n751 & ~n756;
  assign n758 = ~pi022 & n432;
  assign n759 = n662 & n758;
  assign n760 = pi020 & n759;
  assign n761 = n757 & ~n760;
  assign n762 = n745 & n761;
  assign n763 = n722 & n762;
  assign n764 = n417 & n515;
  assign n765 = ~pi009 & n764;
  assign n766 = ~pi009 & pi010;
  assign n767 = pi008 & n707;
  assign n768 = n654 & n767;
  assign n769 = ~pi007 & n768;
  assign n770 = n766 & n769;
  assign n771 = ~n765 & ~n770;
  assign n772 = n702 & ~n771;
  assign n773 = pi018 & ~pi019;
  assign n774 = ~pi021 & n773;
  assign n775 = n725 & n774;
  assign n776 = ~pi011 & ~pi012;
  assign n777 = ~pi013 & n776;
  assign n778 = n510 & n777;
  assign n779 = n346 & n625;
  assign n780 = pi008 & n779;
  assign n781 = ~pi015 & n780;
  assign n782 = n778 & n781;
  assign n783 = ~n775 & ~n782;
  assign n784 = ~pi011 & pi013;
  assign n785 = n508 & n784;
  assign n786 = ~n458 & n705;
  assign n787 = ~n357 & ~n786;
  assign n788 = pi008 & ~n787;
  assign n789 = pi012 & pi014;
  assign n790 = n547 & n789;
  assign n791 = pi011 & n790;
  assign n792 = pi015 & n518;
  assign n793 = n339 & n792;
  assign n794 = ~n791 & ~n793;
  assign n795 = ~n788 & n794;
  assign n796 = ~n785 & n795;
  assign n797 = n700 & ~n796;
  assign n798 = ~n650 & ~n797;
  assign n799 = n783 & n798;
  assign n800 = ~pi011 & pi012;
  assign n801 = n284 & n767;
  assign n802 = ~n458 & n801;
  assign n803 = pi007 & pi010;
  assign n804 = ~pi009 & n803;
  assign n805 = n802 & n804;
  assign n806 = n800 & n805;
  assign n807 = n799 & ~n806;
  assign n808 = ~n772 & n807;
  assign n809 = pi007 & n520;
  assign n810 = n768 & n809;
  assign n811 = n353 & n767;
  assign n812 = ~pi012 & n234;
  assign n813 = pi007 & ~pi009;
  assign n814 = ~pi010 & n813;
  assign n815 = pi011 & n814;
  assign n816 = ~pi011 & n804;
  assign n817 = ~n815 & ~n816;
  assign n818 = n812 & ~n817;
  assign n819 = pi027 & n818;
  assign n820 = n811 & n819;
  assign n821 = pi056 & n269;
  assign n822 = n347 & n821;
  assign n823 = pi025 & n223;
  assign n824 = n822 & n823;
  assign n825 = pi007 & n238;
  assign n826 = ~pi127 & n825;
  assign n827 = pi001 & n269;
  assign n828 = n826 & n827;
  assign n829 = n354 & n828;
  assign n830 = pi000 & n829;
  assign n831 = ~n824 & ~n830;
  assign n832 = ~n820 & n831;
  assign n833 = ~n810 & n832;
  assign n834 = n391 & n482;
  assign n835 = pi020 & n834;
  assign n836 = ~pi023 & n269;
  assign n837 = ~pi017 & n836;
  assign n838 = n835 & n837;
  assign n839 = ~n383 & n838;
  assign n840 = n270 & n373;
  assign n841 = n480 & n840;
  assign n842 = pi023 & n269;
  assign n843 = ~n383 & n842;
  assign n844 = n392 & n482;
  assign n845 = n843 & n844;
  assign n846 = ~n841 & ~n845;
  assign n847 = ~n839 & n846;
  assign n848 = n233 & n654;
  assign n849 = n591 & n848;
  assign n850 = n251 & n462;
  assign n851 = ~n654 & n850;
  assign n852 = ~n849 & ~n851;
  assign n853 = n689 & ~n852;
  assign n854 = ~pi005 & n853;
  assign n855 = n385 & n451;
  assign n856 = n394 & n468;
  assign n857 = n855 & n856;
  assign n858 = pi016 & n857;
  assign n859 = ~n854 & ~n858;
  assign n860 = n847 & n859;
  assign n861 = n833 & n860;
  assign n862 = n808 & n861;
  assign n863 = pi013 & ~pi015;
  assign n864 = n789 & n863;
  assign n865 = ~pi008 & n707;
  assign n866 = n813 & n865;
  assign n867 = ~pi010 & n866;
  assign n868 = n864 & n867;
  assign n869 = n491 & n734;
  assign n870 = pi020 & n869;
  assign n871 = ~pi013 & n579;
  assign n872 = n800 & n871;
  assign n873 = pi007 & n872;
  assign n874 = n865 & n873;
  assign n875 = ~n870 & ~n874;
  assign n876 = ~n868 & n875;
  assign n877 = n862 & n876;
  assign n878 = n763 & n877;
  assign n879 = ~pi090 & ~pi091;
  assign n880 = ~pi092 & n879;
  assign n881 = n446 & n736;
  assign n882 = n880 & n881;
  assign n883 = n677 & n882;
  assign n884 = ~pi093 & n883;
  assign n885 = ~pi094 & n884;
  assign n886 = ~pi095 & n885;
  assign n887 = pi096 & n886;
  assign n888 = pi094 & n884;
  assign n889 = ~n887 & ~n888;
  assign n890 = n802 & n815;
  assign n891 = pi012 & n890;
  assign n892 = n332 & n779;
  assign n893 = n704 & n892;
  assign n894 = n462 & n893;
  assign n895 = n361 & n416;
  assign n896 = n766 & n776;
  assign n897 = n895 & n896;
  assign n898 = ~pi013 & n897;
  assign n899 = ~n894 & ~n898;
  assign n900 = ~n891 & n899;
  assign n901 = n889 & n900;
  assign n902 = n878 & n901;
  assign n903 = ~pi011 & ~pi013;
  assign n904 = ~pi014 & n903;
  assign n905 = n709 & n801;
  assign n906 = pi015 & n905;
  assign n907 = n904 & n906;
  assign n908 = pi010 & ~pi011;
  assign n909 = n708 & n767;
  assign n910 = n654 & n909;
  assign n911 = n908 & n910;
  assign n912 = n284 & n779;
  assign n913 = n871 & n912;
  assign n914 = ~pi008 & pi015;
  assign n915 = ~n339 & ~n914;
  assign n916 = n913 & ~n915;
  assign n917 = ~pi011 & n916;
  assign n918 = ~n911 & ~n917;
  assign n919 = ~n907 & n918;
  assign n920 = n233 & ~n234;
  assign n921 = n867 & ~n920;
  assign n922 = ~pi010 & ~pi011;
  assign n923 = n708 & n865;
  assign n924 = n922 & n923;
  assign n925 = n812 & n924;
  assign n926 = pi011 & ~pi013;
  assign n927 = n510 & n780;
  assign n928 = n812 & n927;
  assign n929 = n926 & n928;
  assign n930 = ~n925 & ~n929;
  assign n931 = ~n921 & n930;
  assign n932 = ~n864 & ~n931;
  assign n933 = n919 & ~n932;
  assign n934 = pi013 & n511;
  assign n935 = n709 & n811;
  assign n936 = pi027 & n935;
  assign n937 = pi014 & n936;
  assign n938 = n934 & n937;
  assign n939 = pi015 & n938;
  assign n940 = ~pi039 & n694;
  assign n941 = n683 & n940;
  assign n942 = ~n631 & ~n941;
  assign n943 = ~n939 & n942;
  assign n944 = n933 & n943;
  assign po05 = ~n902 | ~n944;
  assign n946 = n591 & n659;
  assign n947 = n230 & n408;
  assign n948 = pi023 & n947;
  assign n949 = n267 & n451;
  assign n950 = n948 & n949;
  assign n951 = pi082 & n950;
  assign n952 = n284 & n950;
  assign n953 = ~n951 & ~n952;
  assign n954 = n386 & n626;
  assign n955 = pi057 & n954;
  assign n956 = n953 & ~n955;
  assign n957 = ~pi045 & ~n956;
  assign n958 = pi022 & n773;
  assign n959 = n821 & n958;
  assign n960 = n277 & n959;
  assign n961 = pi023 & n960;
  assign n962 = n353 & n961;
  assign n963 = n277 & n842;
  assign n964 = ~pi036 & n963;
  assign n965 = ~pi035 & n964;
  assign n966 = ~pi022 & n773;
  assign n967 = pi021 & ~pi037;
  assign n968 = n966 & ~n967;
  assign n969 = n965 & n968;
  assign n970 = n277 & n966;
  assign n971 = ~pi035 & pi036;
  assign n972 = n269 & n971;
  assign n973 = n970 & n972;
  assign n974 = ~pi012 & n705;
  assign n975 = n582 & n974;
  assign n976 = ~n973 & ~n975;
  assign n977 = ~n969 & n976;
  assign n978 = ~pi013 & n800;
  assign n979 = n332 & n978;
  assign n980 = ~pi015 & n509;
  assign n981 = n979 & n980;
  assign n982 = pi011 & n418;
  assign n983 = pi012 & n982;
  assign n984 = pi013 & ~pi014;
  assign n985 = pi015 & n984;
  assign n986 = n983 & n985;
  assign n987 = ~n981 & ~n986;
  assign n988 = n419 & ~n458;
  assign n989 = ~n379 & ~n988;
  assign n990 = n666 & n989;
  assign n991 = ~n371 & n990;
  assign n992 = n987 & n991;
  assign n993 = n977 & n992;
  assign n994 = n284 & ~n993;
  assign n995 = ~pi081 & pi083;
  assign n996 = ~pi080 & n995;
  assign n997 = ~pi056 & ~pi082;
  assign n998 = n996 & n997;
  assign n999 = n963 & n998;
  assign n1000 = n353 & n999;
  assign n1001 = ~pi065 & n958;
  assign n1002 = pi021 & n1001;
  assign n1003 = ~n855 & ~n1002;
  assign n1004 = n1000 & ~n1003;
  assign n1005 = n582 & n934;
  assign n1006 = n268 & n625;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n1004 & n1007;
  assign n1009 = ~n994 & n1008;
  assign n1010 = ~n962 & n1009;
  assign n1011 = ~n957 & n1010;
  assign n1012 = ~n946 & n1011;
  assign n1013 = ~n383 & ~n1012;
  assign n1014 = n337 & n347;
  assign n1015 = ~n262 & n1014;
  assign n1016 = ~pi079 & n248;
  assign n1017 = n1014 & ~n1016;
  assign n1018 = ~pi122 & n1017;
  assign n1019 = ~n325 & ~n1018;
  assign n1020 = n332 & n974;
  assign n1021 = pi015 & n580;
  assign n1022 = n1020 & n1021;
  assign n1023 = ~n262 & n1022;
  assign n1024 = ~n365 & ~n1023;
  assign n1025 = n1019 & n1024;
  assign n1026 = ~n1015 & n1025;
  assign n1027 = ~n266 & n1026;
  assign n1028 = n284 & n828;
  assign n1029 = pi000 & n1028;
  assign n1030 = ~n306 & ~n321;
  assign n1031 = ~n400 & n1030;
  assign n1032 = ~n318 & n1031;
  assign n1033 = ~n303 & ~n330;
  assign n1034 = ~n307 & n1033;
  assign n1035 = n1032 & n1034;
  assign n1036 = ~n310 & n1035;
  assign n1037 = ~n355 & n1036;
  assign n1038 = ~n1029 & n1037;
  assign n1039 = ~n302 & ~n1038;
  assign n1040 = n262 & n1035;
  assign n1041 = ~n355 & n1040;
  assign n1042 = n1039 & ~n1041;
  assign n1043 = pi044 & ~n382;
  assign n1044 = pi001 & n494;
  assign n1045 = n825 & n1044;
  assign n1046 = n269 & n1045;
  assign n1047 = n284 & n1046;
  assign n1048 = ~n1043 & n1047;
  assign n1049 = n239 & n309;
  assign n1050 = ~pi001 & n1049;
  assign n1051 = n224 & n1050;
  assign n1052 = ~n1048 & ~n1051;
  assign n1053 = ~n1028 & ~n1049;
  assign n1054 = ~pi122 & ~n1053;
  assign n1055 = n299 & ~n1054;
  assign n1056 = n1052 & n1055;
  assign n1057 = ~n1042 & n1056;
  assign n1058 = n1027 & n1057;
  assign n1059 = ~pi045 & n284;
  assign n1060 = n580 & n778;
  assign n1061 = n1059 & n1060;
  assign n1062 = ~n527 & ~n1061;
  assign n1063 = n274 & n495;
  assign n1064 = n574 & n1063;
  assign n1065 = n251 & n754;
  assign n1066 = n392 & n1065;
  assign n1067 = ~n1064 & ~n1066;
  assign n1068 = ~pi122 & n284;
  assign n1069 = ~n223 & n284;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1067 & ~n1070;
  assign n1072 = n284 & n726;
  assign n1073 = n609 & n1072;
  assign n1074 = n277 & n1073;
  assign n1075 = ~n383 & n1074;
  assign n1076 = ~n1071 & ~n1075;
  assign n1077 = n1062 & n1076;
  assign n1078 = n726 & n948;
  assign n1079 = pi122 & n1078;
  assign n1080 = ~pi122 & n389;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = ~pi002 & n1044;
  assign n1083 = pi003 & ~pi007;
  assign n1084 = n1082 & n1083;
  assign n1085 = pi004 & ~pi006;
  assign n1086 = ~n250 & ~n1085;
  assign n1087 = n1084 & n1086;
  assign n1088 = ~n383 & n1087;
  assign n1089 = ~n234 & ~n515;
  assign n1090 = n333 & n461;
  assign n1091 = n229 & n1090;
  assign n1092 = ~n1089 & n1091;
  assign n1093 = ~n1088 & ~n1092;
  assign n1094 = n408 & n476;
  assign n1095 = n551 & n1094;
  assign n1096 = n270 & n375;
  assign n1097 = pi020 & n391;
  assign n1098 = n432 & n1097;
  assign n1099 = n1096 & n1098;
  assign n1100 = n408 & n432;
  assign n1101 = n966 & n1100;
  assign n1102 = ~n1099 & ~n1101;
  assign n1103 = ~n1095 & n1102;
  assign n1104 = n1093 & n1103;
  assign n1105 = n1081 & n1104;
  assign n1106 = n251 & n661;
  assign n1107 = n881 & n1106;
  assign n1108 = ~pi020 & n276;
  assign n1109 = ~pi017 & n1108;
  assign n1110 = n387 & n540;
  assign n1111 = n1109 & n1110;
  assign n1112 = pi022 & n1111;
  assign n1113 = pi019 & n1112;
  assign n1114 = ~n1107 & ~n1113;
  assign n1115 = ~n1070 & ~n1114;
  assign n1116 = ~n342 & ~n399;
  assign n1117 = n225 & n560;
  assign n1118 = ~n1116 & n1117;
  assign n1119 = ~n383 & n1118;
  assign n1120 = ~n1115 & ~n1119;
  assign n1121 = n1105 & n1120;
  assign n1122 = n1077 & n1121;
  assign n1123 = n251 & n472;
  assign n1124 = n451 & n1123;
  assign n1125 = n469 & n1124;
  assign n1126 = pi017 & n391;
  assign n1127 = n270 & n1126;
  assign n1128 = n387 & n407;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = ~n626 & n1129;
  assign n1131 = n1123 & ~n1130;
  assign n1132 = ~n1125 & ~n1131;
  assign n1133 = ~n383 & ~n1132;
  assign n1134 = ~pi022 & n1111;
  assign n1135 = ~pi023 & n591;
  assign n1136 = n491 & n1135;
  assign n1137 = ~pi005 & n1136;
  assign n1138 = n392 & n1137;
  assign n1139 = ~n1134 & ~n1138;
  assign n1140 = n229 & n1045;
  assign n1141 = n250 & n1063;
  assign n1142 = n346 & n1082;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n497 & n1143;
  assign n1145 = ~n1140 & n1144;
  assign n1146 = n1139 & n1145;
  assign n1147 = ~n383 & ~n1146;
  assign n1148 = ~n614 & ~n1147;
  assign n1149 = pi019 & n374;
  assign n1150 = n408 & n1149;
  assign n1151 = pi018 & n471;
  assign n1152 = n375 & n1151;
  assign n1153 = pi019 & n451;
  assign n1154 = n471 & n1153;
  assign n1155 = ~n1152 & ~n1154;
  assign n1156 = ~n1150 & n1155;
  assign n1157 = n551 & ~n1156;
  assign n1158 = n230 & n461;
  assign n1159 = n235 & n1158;
  assign n1160 = ~n1157 & ~n1159;
  assign n1161 = n1148 & n1160;
  assign n1162 = ~n1133 & n1161;
  assign n1163 = n1122 & n1162;
  assign n1164 = pi055 & pi056;
  assign n1165 = pi122 & n1164;
  assign n1166 = n284 & ~n1165;
  assign n1167 = pi046 & n244;
  assign n1168 = n251 & n1167;
  assign n1169 = n1166 & n1168;
  assign n1170 = n247 & n248;
  assign n1171 = ~pi112 & n533;
  assign n1172 = n244 & n1171;
  assign n1173 = ~n1166 & ~n1172;
  assign n1174 = n1170 & ~n1173;
  assign n1175 = ~n1169 & ~n1174;
  assign n1176 = n254 & n1016;
  assign n1177 = ~n616 & ~n1176;
  assign n1178 = n1166 & ~n1177;
  assign n1179 = n1175 & ~n1178;
  assign n1180 = ~n281 & n1179;
  assign n1181 = n538 & n1180;
  assign n1182 = ~pi006 & n598;
  assign n1183 = ~n383 & n581;
  assign n1184 = pi011 & n547;
  assign n1185 = ~pi011 & n863;
  assign n1186 = ~pi011 & pi015;
  assign n1187 = n462 & ~n1186;
  assign n1188 = ~n1185 & ~n1187;
  assign n1189 = ~n1184 & n1188;
  assign n1190 = n1183 & ~n1189;
  assign n1191 = ~n1182 & ~n1190;
  assign n1192 = n489 & n1191;
  assign n1193 = n384 & n392;
  assign n1194 = ~pi020 & pi022;
  assign n1195 = n1193 & ~n1194;
  assign n1196 = n1153 & n1195;
  assign n1197 = n467 & n553;
  assign n1198 = n948 & n1197;
  assign n1199 = ~pi001 & n460;
  assign n1200 = n345 & n1199;
  assign n1201 = pi019 & n387;
  assign n1202 = n343 & n369;
  assign n1203 = n1201 & n1202;
  assign n1204 = ~n1200 & ~n1203;
  assign n1205 = ~n1198 & n1204;
  assign n1206 = ~n1196 & n1205;
  assign n1207 = ~pi045 & ~n1206;
  assign n1208 = ~pi015 & n418;
  assign n1209 = ~pi012 & n904;
  assign n1210 = n1208 & n1209;
  assign n1211 = ~pi100 & n1210;
  assign n1212 = n1014 & n1068;
  assign n1213 = n1016 & n1212;
  assign n1214 = ~n287 & ~n1213;
  assign n1215 = ~n1211 & n1214;
  assign n1216 = ~n491 & ~n678;
  assign n1217 = ~pi045 & n570;
  assign n1218 = ~n1216 & n1217;
  assign n1219 = n1215 & ~n1218;
  assign n1220 = ~n1207 & n1219;
  assign n1221 = n353 & ~n522;
  assign n1222 = n524 & n1221;
  assign n1223 = ~pi027 & n1222;
  assign n1224 = ~pi014 & n801;
  assign n1225 = pi012 & n814;
  assign n1226 = n1224 & n1225;
  assign n1227 = n1185 & n1226;
  assign n1228 = n458 & n982;
  assign n1229 = pi012 & n1228;
  assign n1230 = ~pi122 & n1229;
  assign n1231 = ~n1227 & ~n1230;
  assign n1232 = ~n1223 & n1231;
  assign n1233 = n557 & n948;
  assign po67 = n272 & n1126;
  assign n1235 = n407 & n837;
  assign n1236 = n1096 & n1235;
  assign n1237 = ~po67 & ~n1236;
  assign n1238 = ~n1233 & n1237;
  assign n1239 = n758 & n840;
  assign n1240 = ~n759 & ~n1239;
  assign n1241 = ~pi015 & n463;
  assign n1242 = n230 & n1241;
  assign n1243 = pi006 & ~pi007;
  assign n1244 = n345 & n1243;
  assign n1245 = n1082 & n1244;
  assign n1246 = ~n383 & n1245;
  assign n1247 = ~n1242 & ~n1246;
  assign n1248 = n284 & n473;
  assign n1249 = n408 & n1248;
  assign n1250 = n443 & n1249;
  assign n1251 = n1247 & ~n1250;
  assign n1252 = n1240 & n1251;
  assign n1253 = n1238 & n1252;
  assign n1254 = n1232 & n1253;
  assign n1255 = n1220 & n1254;
  assign n1256 = n1192 & n1255;
  assign n1257 = n1181 & n1256;
  assign n1258 = n334 & n416;
  assign n1259 = n579 & n1258;
  assign n1260 = n914 & n1259;
  assign n1261 = ~pi007 & n579;
  assign n1262 = n767 & n1261;
  assign n1263 = pi014 & n1262;
  assign n1264 = n776 & n1263;
  assign n1265 = ~n284 & n343;
  assign n1266 = pi019 & n277;
  assign n1267 = n270 & n1266;
  assign n1268 = n433 & n1267;
  assign n1269 = ~n593 & ~n1268;
  assign n1270 = n1265 & ~n1269;
  assign n1271 = n235 & n982;
  assign n1272 = ~n284 & n1271;
  assign n1273 = ~n1270 & ~n1272;
  assign n1274 = ~n1264 & n1273;
  assign n1275 = ~n1260 & n1274;
  assign n1276 = n469 & n609;
  assign n1277 = ~n383 & n1276;
  assign n1278 = n374 & n472;
  assign n1279 = ~n1197 & ~n1278;
  assign n1280 = n1277 & ~n1279;
  assign n1281 = n392 & n551;
  assign n1282 = n678 & n1281;
  assign n1283 = n392 & n1197;
  assign n1284 = n551 & n1283;
  assign n1285 = n373 & n551;
  assign n1286 = n774 & n1285;
  assign n1287 = ~n1284 & ~n1286;
  assign n1288 = ~n1282 & n1287;
  assign n1289 = ~n1280 & n1288;
  assign n1290 = ~n383 & n418;
  assign n1291 = n512 & n1290;
  assign n1292 = n423 & n659;
  assign n1293 = n443 & n1267;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n1291 & n1294;
  assign n1296 = n1289 & n1295;
  assign n1297 = n1275 & n1296;
  assign n1298 = n269 & n474;
  assign n1299 = n225 & n1044;
  assign n1300 = pi007 & n1299;
  assign n1301 = n230 & n1300;
  assign n1302 = n473 & n1276;
  assign n1303 = n609 & n1109;
  assign n1304 = pi022 & n387;
  assign n1305 = n1303 & n1304;
  assign n1306 = n269 & n1084;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1302 & n1307;
  assign n1309 = ~n1301 & n1308;
  assign n1310 = ~n1043 & ~n1309;
  assign n1311 = ~n1298 & ~n1310;
  assign n1312 = n269 & n291;
  assign n1313 = n354 & n1312;
  assign n1314 = ~n1164 & n1313;
  assign n1315 = pi122 & ~n1164;
  assign n1316 = n284 & n1315;
  assign n1317 = n319 & n320;
  assign n1318 = n1316 & n1317;
  assign n1319 = ~n1314 & ~n1318;
  assign n1320 = n278 & n959;
  assign n1321 = ~n1070 & n1320;
  assign n1322 = n1319 & ~n1321;
  assign n1323 = pi025 & n404;
  assign n1324 = ~pi024 & n1323;
  assign n1325 = ~n282 & ~n1324;
  assign n1326 = n1020 & ~n1325;
  assign n1327 = n769 & n1326;
  assign n1328 = n517 & n979;
  assign n1329 = n284 & n1328;
  assign n1330 = ~n1327 & ~n1329;
  assign n1331 = ~n383 & n947;
  assign n1332 = n376 & n1331;
  assign n1333 = n1330 & ~n1332;
  assign n1334 = pi004 & n291;
  assign n1335 = n308 & n1334;
  assign n1336 = ~n637 & ~n1335;
  assign n1337 = ~n1312 & n1336;
  assign n1338 = n292 & n343;
  assign n1339 = n1337 & ~n1338;
  assign n1340 = n1069 & ~n1339;
  assign n1341 = ~pi007 & n425;
  assign n1342 = n317 & n1341;
  assign n1343 = pi061 & n1342;
  assign n1344 = ~n1165 & n1343;
  assign n1345 = ~pi061 & n1342;
  assign n1346 = pi027 & n618;
  assign n1347 = n1312 & n1346;
  assign n1348 = ~n223 & n1347;
  assign n1349 = ~n1345 & ~n1348;
  assign n1350 = ~n1344 & n1349;
  assign n1351 = ~n1340 & n1350;
  assign n1352 = n1333 & n1351;
  assign n1353 = n1322 & n1352;
  assign n1354 = n1311 & n1353;
  assign n1355 = n1297 & n1354;
  assign n1356 = n230 & n573;
  assign n1357 = ~n284 & n1356;
  assign n1358 = n411 & n1265;
  assign n1359 = n267 & n270;
  assign n1360 = n284 & n677;
  assign n1361 = n1359 & n1360;
  assign n1362 = ~n1358 & ~n1361;
  assign n1363 = pi023 & ~n1362;
  assign n1364 = pi088 & ~pi117;
  assign n1365 = n533 & n1364;
  assign n1366 = n625 & n1365;
  assign n1367 = ~n1363 & ~n1366;
  assign n1368 = ~n1357 & n1367;
  assign n1369 = pi013 & n896;
  assign n1370 = n339 & n1369;
  assign n1371 = n416 & n1370;
  assign n1372 = pi125 & ~pi126;
  assign n1373 = n353 & n1372;
  assign n1374 = ~n1371 & ~n1373;
  assign n1375 = ~n596 & n1374;
  assign n1376 = ~n579 & n702;
  assign n1377 = ~n766 & n1376;
  assign n1378 = n517 & n1377;
  assign n1379 = n343 & n689;
  assign n1380 = ~n333 & n1379;
  assign n1381 = ~n1378 & ~n1380;
  assign n1382 = n1375 & n1381;
  assign n1383 = ~pi018 & n472;
  assign n1384 = n485 & n1383;
  assign n1385 = n392 & n855;
  assign n1386 = n483 & n1385;
  assign n1387 = pi020 & n1386;
  assign n1388 = ~n1384 & ~n1387;
  assign n1389 = n228 & n1244;
  assign n1390 = n684 & n1389;
  assign n1391 = n647 & n790;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = n234 & n974;
  assign n1394 = n418 & n1393;
  assign n1395 = n1392 & ~n1394;
  assign n1396 = n368 & n676;
  assign n1397 = n353 & n1396;
  assign n1398 = n754 & n1397;
  assign n1399 = n872 & n980;
  assign n1400 = n414 & n495;
  assign n1401 = n337 & n1400;
  assign n1402 = ~n1399 & ~n1401;
  assign n1403 = ~n1398 & n1402;
  assign n1404 = n1395 & n1403;
  assign n1405 = n1388 & n1404;
  assign n1406 = n1382 & n1405;
  assign n1407 = n1368 & n1406;
  assign n1408 = ~pi020 & pi021;
  assign n1409 = pi023 & n736;
  assign n1410 = ~pi022 & n1409;
  assign n1411 = n1408 & n1410;
  assign n1412 = n661 & n1411;
  assign n1413 = n269 & n1412;
  assign n1414 = ~pi021 & n736;
  assign n1415 = n369 & n1414;
  assign n1416 = pi022 & n836;
  assign n1417 = n1415 & n1416;
  assign n1418 = ~n1228 & ~n1417;
  assign n1419 = pi047 & n359;
  assign n1420 = pi113 & n1419;
  assign n1421 = n362 & n1420;
  assign n1422 = n354 & n1421;
  assign n1423 = n1418 & ~n1422;
  assign n1424 = ~n1413 & n1423;
  assign n1425 = n224 & ~n1424;
  assign n1426 = n284 & n483;
  assign n1427 = ~n627 & ~n1268;
  assign n1428 = n226 & n592;
  assign n1429 = pi003 & n1428;
  assign n1430 = ~n411 & ~n1429;
  assign n1431 = n1427 & n1430;
  assign n1432 = n1426 & ~n1431;
  assign n1433 = ~n645 & ~n1356;
  assign n1434 = ~n1070 & ~n1433;
  assign n1435 = ~n1432 & ~n1434;
  assign n1436 = ~n1425 & n1435;
  assign n1437 = n651 & ~n1070;
  assign n1438 = n1359 & n1396;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~pi023 & n737;
  assign n1441 = n1396 & n1440;
  assign n1442 = pi021 & n1441;
  assign n1443 = n224 & n435;
  assign n1444 = ~n737 & ~n752;
  assign n1445 = n609 & ~n1444;
  assign n1446 = n1443 & n1445;
  assign n1447 = n678 & n836;
  assign n1448 = n1443 & n1447;
  assign n1449 = ~n1446 & ~n1448;
  assign n1450 = ~n1442 & n1449;
  assign n1451 = n271 & n472;
  assign n1452 = n391 & n1451;
  assign n1453 = ~n273 & n1452;
  assign n1454 = n895 & n979;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = n361 & n1259;
  assign n1457 = n1455 & ~n1456;
  assign n1458 = n473 & n570;
  assign n1459 = n273 & n676;
  assign n1460 = n754 & n1459;
  assign n1461 = ~n1458 & ~n1460;
  assign n1462 = n1457 & n1461;
  assign n1463 = n1450 & n1462;
  assign n1464 = ~n648 & ~n792;
  assign n1465 = n647 & ~n1464;
  assign n1466 = n414 & n685;
  assign n1467 = ~n383 & n1466;
  assign n1468 = ~n1465 & ~n1467;
  assign n1469 = ~pi021 & n1440;
  assign n1470 = n435 & n1469;
  assign n1471 = n1426 & n1470;
  assign n1472 = n1468 & ~n1471;
  assign n1473 = n461 & n518;
  assign n1474 = ~pi014 & n1473;
  assign n1475 = n346 & n1474;
  assign n1476 = n1069 & n1475;
  assign n1477 = ~pi013 & n789;
  assign n1478 = pi011 & n1477;
  assign n1479 = pi008 & n892;
  assign n1480 = n1478 & n1479;
  assign n1481 = pi012 & n546;
  assign n1482 = n654 & n1481;
  assign n1483 = n333 & n1089;
  assign n1484 = n1158 & n1483;
  assign n1485 = ~n1482 & ~n1484;
  assign n1486 = ~n1480 & n1485;
  assign n1487 = ~n1476 & n1486;
  assign n1488 = n1472 & n1487;
  assign n1489 = n1463 & n1488;
  assign n1490 = n1439 & n1489;
  assign n1491 = n1436 & n1490;
  assign n1492 = n1407 & n1491;
  assign n1493 = n1355 & n1492;
  assign n1494 = n1257 & n1493;
  assign n1495 = n1163 & n1494;
  assign n1496 = n1058 & n1495;
  assign n1497 = ~pi096 & n886;
  assign n1498 = pi023 & n385;
  assign n1499 = pi017 & ~pi018;
  assign n1500 = n1498 & n1499;
  assign n1501 = n676 & n1500;
  assign n1502 = n880 & n1501;
  assign n1503 = ~pi021 & n1502;
  assign n1504 = n882 & n1396;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = ~n1497 & n1505;
  assign n1507 = ~pi097 & ~pi098;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = pi093 & n883;
  assign n1510 = pi095 & n885;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n880 & n1501;
  assign n1513 = n1511 & ~n1512;
  assign n1514 = n889 & n1513;
  assign n1515 = ~n1508 & n1514;
  assign n1516 = n423 & n1341;
  assign n1517 = ~n576 & ~n1516;
  assign n1518 = pi039 & n575;
  assign n1519 = n1517 & ~n1518;
  assign n1520 = n1515 & n1519;
  assign n1521 = n573 & n1426;
  assign n1522 = ~n810 & ~n1521;
  assign n1523 = ~n397 & n1522;
  assign n1524 = n1520 & n1523;
  assign n1525 = n408 & n752;
  assign n1526 = ~pi022 & n1525;
  assign n1527 = n482 & n1109;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = n443 & ~n1528;
  assign n1530 = n1524 & ~n1529;
  assign n1531 = n437 & n609;
  assign n1532 = ~pi122 & n1531;
  assign n1533 = n1201 & n1303;
  assign n1534 = n1110 & n1266;
  assign n1535 = pi022 & n1534;
  assign n1536 = ~pi022 & n387;
  assign n1537 = n251 & n1266;
  assign n1538 = n1536 & n1537;
  assign n1539 = ~n1535 & ~n1538;
  assign n1540 = ~n1533 & n1539;
  assign n1541 = ~pi122 & ~n1540;
  assign n1542 = ~pi122 & n609;
  assign n1543 = n1097 & n1201;
  assign n1544 = n1542 & n1543;
  assign n1545 = ~pi122 & n748;
  assign n1546 = n1303 & n1545;
  assign n1547 = pi005 & pi006;
  assign n1548 = n1300 & n1547;
  assign n1549 = ~pi122 & n1548;
  assign n1550 = n269 & n560;
  assign n1551 = ~pi122 & n1550;
  assign n1552 = pi002 & n494;
  assign n1553 = n827 & n1552;
  assign n1554 = ~pi122 & n1553;
  assign n1555 = ~n1551 & ~n1554;
  assign n1556 = ~n1549 & n1555;
  assign n1557 = ~n1546 & n1556;
  assign n1558 = ~n1544 & n1557;
  assign n1559 = ~n1541 & n1558;
  assign n1560 = ~n1532 & n1559;
  assign n1561 = ~pi023 & n1201;
  assign n1562 = ~pi022 & n1561;
  assign n1563 = n1106 & n1562;
  assign n1564 = ~n1534 & ~n1563;
  assign n1565 = n632 & n1201;
  assign n1566 = n1564 & ~n1565;
  assign n1567 = n1108 & n1137;
  assign n1568 = n271 & n436;
  assign n1569 = ~pi003 & n1550;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1567 & n1570;
  assign n1572 = n1566 & n1571;
  assign n1573 = n224 & ~n1572;
  assign n1574 = pi004 & n1300;
  assign n1575 = n224 & n1574;
  assign n1576 = ~pi005 & n1574;
  assign n1577 = ~pi122 & n1576;
  assign n1578 = ~n1575 & ~n1577;
  assign n1579 = n434 & n834;
  assign n1580 = n251 & n1579;
  assign n1581 = pi017 & n834;
  assign n1582 = n541 & n1581;
  assign n1583 = ~n1580 & ~n1582;
  assign n1584 = ~pi122 & ~n1583;
  assign n1585 = n224 & n251;
  assign n1586 = n1581 & n1585;
  assign n1587 = ~n1584 & ~n1586;
  assign n1588 = pi003 & n1553;
  assign n1589 = n224 & n1588;
  assign n1590 = n1587 & ~n1589;
  assign n1591 = n1578 & n1590;
  assign n1592 = ~n1573 & n1591;
  assign n1593 = n1560 & n1592;
  assign n1594 = n471 & n569;
  assign n1595 = ~n673 & ~n1594;
  assign n1596 = ~n410 & n1595;
  assign n1597 = n480 & ~n1596;
  assign n1598 = pi021 & pi022;
  assign n1599 = pi019 & n1598;
  assign n1600 = n392 & n1599;
  assign n1601 = ~n749 & n1600;
  assign n1602 = n391 & n749;
  assign n1603 = n557 & n1602;
  assign n1604 = ~n558 & ~n1603;
  assign n1605 = ~n1601 & n1604;
  assign n1606 = n480 & ~n1605;
  assign n1607 = n373 & n480;
  assign n1608 = ~n270 & ~n557;
  assign n1609 = n1607 & ~n1608;
  assign n1610 = pi018 & pi019;
  assign n1611 = n1607 & n1610;
  assign n1612 = ~n1598 & n1611;
  assign n1613 = ~n1609 & ~n1612;
  assign n1614 = ~n1606 & n1613;
  assign n1615 = ~n1597 & n1614;
  assign n1616 = ~n493 & n1615;
  assign n1617 = n1316 & n1421;
  assign n1618 = n284 & n343;
  assign n1619 = ~pi019 & n374;
  assign n1620 = n433 & n1619;
  assign n1621 = n1364 & n1620;
  assign n1622 = n1618 & n1621;
  assign n1623 = n373 & n1622;
  assign n1624 = ~n1617 & ~n1623;
  assign n1625 = n284 & n392;
  assign n1626 = n1536 & n1625;
  assign n1627 = n588 & n1626;
  assign n1628 = n1624 & ~n1627;
  assign n1629 = n1616 & n1628;
  assign n1630 = pi001 & pi003;
  assign n1631 = n1552 & n1630;
  assign n1632 = ~n383 & n1631;
  assign n1633 = ~n1116 & n1632;
  assign n1634 = n1629 & ~n1633;
  assign n1635 = n1593 & n1634;
  assign n1636 = n1068 & n1317;
  assign n1637 = n386 & n672;
  assign n1638 = n224 & n1637;
  assign n1639 = n736 & n947;
  assign n1640 = n224 & n1639;
  assign n1641 = ~n1598 & n1640;
  assign n1642 = ~n1638 & ~n1641;
  assign n1643 = n391 & n1197;
  assign n1644 = n588 & n1643;
  assign n1645 = ~n635 & ~n1644;
  assign n1646 = n452 & n678;
  assign n1647 = n588 & n1646;
  assign n1648 = n551 & n1415;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = n1645 & n1649;
  assign n1651 = n542 & n748;
  assign n1652 = ~n383 & n1651;
  assign n1653 = n546 & n812;
  assign n1654 = ~pi014 & n229;
  assign n1655 = ~n230 & ~n1654;
  assign n1656 = n1473 & ~n1655;
  assign n1657 = ~n1653 & ~n1656;
  assign n1658 = ~n1652 & n1657;
  assign n1659 = n550 & n1658;
  assign n1660 = n1650 & n1659;
  assign n1661 = ~pi122 & n1639;
  assign n1662 = n1660 & ~n1661;
  assign n1663 = n1642 & n1662;
  assign n1664 = pi007 & n425;
  assign n1665 = n1109 & n1359;
  assign n1666 = ~n500 & ~n1665;
  assign n1667 = ~pi019 & n626;
  assign n1668 = n1666 & ~n1667;
  assign n1669 = ~n1664 & n1668;
  assign n1670 = n435 & n1197;
  assign n1671 = n1669 & ~n1670;
  assign n1672 = n483 & ~n1671;
  assign n1673 = n251 & n1152;
  assign n1674 = n586 & n1673;
  assign n1675 = n452 & n748;
  assign n1676 = n540 & n1675;
  assign n1677 = ~n383 & n1676;
  assign n1678 = n540 & n844;
  assign n1679 = n342 & n1045;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = ~n383 & ~n1680;
  assign n1682 = ~n1677 & ~n1681;
  assign n1683 = ~n1674 & n1682;
  assign n1684 = n1409 & n1459;
  assign n1685 = n1683 & ~n1684;
  assign n1686 = ~n572 & n1685;
  assign n1687 = ~n1672 & n1686;
  assign n1688 = n1663 & n1687;
  assign n1689 = ~n1636 & n1688;
  assign n1690 = n1635 & n1689;
  assign n1691 = n1530 & n1690;
  assign n1692 = n1496 & n1691;
  assign po06 = n1013 | ~n1692;
  assign n1694 = n224 & n1568;
  assign n1695 = n224 & n1567;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = n224 & n1569;
  assign n1698 = ~pi002 & n1697;
  assign n1699 = n1696 & ~n1698;
  assign n1700 = n333 & n1263;
  assign n1701 = pi015 & n1700;
  assign n1702 = ~pi011 & n1701;
  assign n1703 = n508 & n779;
  assign n1704 = n360 & n1703;
  assign n1705 = n542 & n1536;
  assign n1706 = n354 & n1705;
  assign n1707 = n269 & n463;
  assign n1708 = ~n515 & n1707;
  assign n1709 = ~n1706 & ~n1708;
  assign n1710 = ~n1704 & n1709;
  assign n1711 = ~n1702 & n1710;
  assign n1712 = n1100 & n1201;
  assign n1713 = ~pi022 & n1712;
  assign n1714 = ~n1674 & ~n1713;
  assign n1715 = n1711 & n1714;
  assign n1716 = n1699 & n1715;
  assign n1717 = pi019 & n760;
  assign n1718 = ~pi008 & n458;
  assign n1719 = n979 & n1718;
  assign n1720 = n416 & n1719;
  assign n1721 = ~n829 & ~n1720;
  assign n1722 = ~n1717 & n1721;
  assign n1723 = pi039 & n230;
  assign n1724 = n284 & n496;
  assign n1725 = n1723 & n1724;
  assign n1726 = n1276 & n1278;
  assign n1727 = n224 & n1726;
  assign n1728 = ~pi039 & n284;
  assign n1729 = n231 & n1728;
  assign n1730 = n495 & n1729;
  assign n1731 = ~n1727 & ~n1730;
  assign n1732 = ~n1725 & n1731;
  assign n1733 = n1722 & n1732;
  assign n1734 = ~pi014 & n1262;
  assign n1735 = ~pi015 & n358;
  assign n1736 = ~n903 & ~n1735;
  assign n1737 = n1734 & ~n1736;
  assign n1738 = n1733 & ~n1737;
  assign n1739 = pi108 & ~pi109;
  assign n1740 = n317 & n1045;
  assign n1741 = pi021 & n472;
  assign n1742 = n540 & n1741;
  assign n1743 = n1151 & n1742;
  assign n1744 = ~n1740 & ~n1743;
  assign n1745 = n284 & ~n1744;
  assign n1746 = pi045 & n1745;
  assign n1747 = n1739 & n1746;
  assign n1748 = pi009 & n780;
  assign n1749 = n462 & n1748;
  assign n1750 = ~pi014 & n908;
  assign n1751 = n1749 & ~n1750;
  assign n1752 = ~n1747 & ~n1751;
  assign n1753 = n1738 & n1752;
  assign n1754 = n1716 & n1753;
  assign n1755 = n491 & n570;
  assign n1756 = pi023 & n1383;
  assign n1757 = n747 & n1756;
  assign n1758 = ~n1755 & ~n1757;
  assign n1759 = n570 & n1536;
  assign n1760 = n354 & n1112;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = ~n1203 & n1761;
  assign n1763 = n1758 & n1762;
  assign n1764 = n373 & n552;
  assign n1765 = ~n1581 & ~n1764;
  assign n1766 = n540 & ~n1765;
  assign n1767 = n541 & n1643;
  assign n1768 = pi017 & n1767;
  assign n1769 = n238 & n1044;
  assign n1770 = ~n316 & n1769;
  assign n1771 = ~n1006 & ~n1770;
  assign n1772 = pi006 & ~n1771;
  assign n1773 = ~n1768 & ~n1772;
  assign n1774 = ~n1766 & n1773;
  assign n1775 = ~n1141 & n1774;
  assign n1776 = ~n383 & ~n1775;
  assign n1777 = pi020 & ~pi021;
  assign n1778 = n1126 & n1777;
  assign n1779 = n476 & n1778;
  assign n1780 = n432 & n1779;
  assign n1781 = ~n1776 & ~n1780;
  assign n1782 = n1763 & n1781;
  assign n1783 = n1754 & n1782;
  assign n1784 = ~n482 & ~n1561;
  assign n1785 = ~pi020 & n747;
  assign n1786 = n284 & n1785;
  assign n1787 = ~n1784 & n1786;
  assign n1788 = n284 & n341;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = n904 & n927;
  assign n1791 = ~pi010 & n1718;
  assign n1792 = n358 & n1791;
  assign n1793 = n912 & n1792;
  assign n1794 = ~pi009 & n1793;
  assign n1795 = ~n1790 & ~n1794;
  assign n1796 = n899 & n1795;
  assign n1797 = n975 & ~n1070;
  assign n1798 = n1796 & ~n1797;
  assign n1799 = n1789 & n1798;
  assign n1800 = ~pi023 & n627;
  assign n1801 = n1426 & n1800;
  assign n1802 = n1285 & n1536;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = n1527 & n1542;
  assign n1805 = ~n1250 & ~n1804;
  assign n1806 = n758 & n1414;
  assign n1807 = n661 & n1806;
  assign n1808 = n1805 & ~n1807;
  assign n1809 = ~n1239 & n1808;
  assign n1810 = n1803 & n1809;
  assign n1811 = n1799 & n1810;
  assign n1812 = n1100 & n1197;
  assign n1813 = n505 & ~n1812;
  assign n1814 = ~pi023 & ~n1813;
  assign n1815 = n334 & n768;
  assign n1816 = n510 & n1815;
  assign n1817 = ~pi007 & n1816;
  assign n1818 = n1542 & n1741;
  assign n1819 = n469 & n1818;
  assign n1820 = ~n1532 & ~n1546;
  assign n1821 = ~n1819 & n1820;
  assign n1822 = ~n1817 & n1821;
  assign n1823 = ~n1814 & n1822;
  assign n1824 = n1811 & n1823;
  assign n1825 = n1126 & n1153;
  assign n1826 = pi020 & n1825;
  assign n1827 = n471 & n1201;
  assign n1828 = ~n835 & ~n1827;
  assign n1829 = ~n1826 & n1828;
  assign n1830 = n551 & ~n1829;
  assign n1831 = n337 & n1474;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n251 & n461;
  assign n1834 = ~pi012 & ~pi014;
  assign n1835 = n547 & n1834;
  assign n1836 = n1833 & n1835;
  assign n1837 = ~n1521 & ~n1836;
  assign n1838 = n777 & n892;
  assign n1839 = ~n458 & n1838;
  assign n1840 = n654 & n1090;
  assign n1841 = n337 & n1840;
  assign n1842 = ~n1839 & ~n1841;
  assign n1843 = n1837 & n1842;
  assign n1844 = n1832 & n1843;
  assign n1845 = pi027 & n1222;
  assign n1846 = pi003 & n494;
  assign n1847 = ~pi001 & n1846;
  assign n1848 = ~pi002 & n1847;
  assign n1849 = ~n229 & ~n345;
  assign n1850 = n424 & ~n1849;
  assign n1851 = n1848 & ~n1850;
  assign n1852 = ~n1446 & ~n1851;
  assign n1853 = ~n1845 & n1852;
  assign n1854 = n423 & n496;
  assign n1855 = ~n1391 & ~n1854;
  assign n1856 = n471 & n1073;
  assign n1857 = n597 & n1084;
  assign n1858 = n619 & n1372;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~n1856 & n1859;
  assign n1861 = n1855 & n1860;
  assign n1862 = ~n383 & n1123;
  assign n1863 = n484 & n1862;
  assign n1864 = pi022 & n1281;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = n270 & ~n1865;
  assign n1867 = n1861 & ~n1866;
  assign n1868 = n483 & n1665;
  assign n1869 = n269 & n284;
  assign n1870 = n234 & n1869;
  assign n1871 = n1473 & n1870;
  assign n1872 = n684 & n1833;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = ~n1868 & n1873;
  assign n1875 = ~pi012 & n458;
  assign n1876 = n705 & n1875;
  assign n1877 = n1479 & n1876;
  assign n1878 = pi019 & n270;
  assign n1879 = n1396 & n1878;
  assign n1880 = ~n1877 & ~n1879;
  assign n1881 = n289 & ~n383;
  assign n1882 = n317 & n1881;
  assign n1883 = n274 & n1882;
  assign n1884 = ~pi127 & n1883;
  assign n1885 = ~pi000 & n1884;
  assign n1886 = n1880 & ~n1885;
  assign n1887 = n1874 & n1886;
  assign n1888 = n1867 & n1887;
  assign n1889 = n508 & n707;
  assign n1890 = n863 & n896;
  assign n1891 = n1889 & n1890;
  assign n1892 = ~pi007 & n1891;
  assign n1893 = n519 & n579;
  assign n1894 = n361 & n1893;
  assign n1895 = n779 & n1894;
  assign n1896 = pi054 & n1895;
  assign n1897 = n284 & n1895;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1892 & n1898;
  assign n1900 = n892 & n1718;
  assign n1901 = n705 & n1900;
  assign n1902 = n518 & n1479;
  assign n1903 = ~n458 & n1902;
  assign n1904 = n776 & n1479;
  assign n1905 = n458 & n1904;
  assign n1906 = ~n1903 & ~n1905;
  assign n1907 = ~n1901 & n1906;
  assign n1908 = n1899 & n1907;
  assign n1909 = n1888 & n1908;
  assign n1910 = n1853 & n1909;
  assign n1911 = n1844 & n1910;
  assign n1912 = n1824 & n1911;
  assign n1913 = n1783 & n1912;
  assign n1914 = ~pi045 & ~pi122;
  assign n1915 = n1739 & n1914;
  assign n1916 = n1745 & n1915;
  assign n1917 = n317 & n1063;
  assign n1918 = ~pi039 & n1917;
  assign n1919 = pi039 & n1917;
  assign n1920 = ~pi049 & n1919;
  assign n1921 = ~n1918 & ~n1920;
  assign n1922 = pi049 & n1919;
  assign n1923 = ~pi051 & n1922;
  assign n1924 = n1921 & ~n1923;
  assign n1925 = n1739 & n1923;
  assign n1926 = ~pi122 & ~n1925;
  assign n1927 = ~n1924 & ~n1926;
  assign n1928 = n484 & n1124;
  assign n1929 = n1921 & ~n1928;
  assign n1930 = ~pi045 & pi122;
  assign n1931 = n1739 & ~n1930;
  assign n1932 = ~n1929 & n1931;
  assign n1933 = ~n1927 & ~n1932;
  assign n1934 = ~n1916 & n1933;
  assign n1935 = ~pi108 & ~pi122;
  assign n1936 = ~pi122 & ~n1935;
  assign n1937 = ~n1745 & ~n1928;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = n686 & n848;
  assign n1940 = ~n751 & ~n1200;
  assign n1941 = n1917 & n1935;
  assign n1942 = n376 & n471;
  assign n1943 = n551 & n1942;
  assign n1944 = ~n1941 & ~n1943;
  assign n1945 = n1940 & n1944;
  assign n1946 = ~n1939 & n1945;
  assign n1947 = ~n1938 & n1946;
  assign n1948 = n1934 & n1947;
  assign n1949 = n337 & n689;
  assign n1950 = n229 & n689;
  assign n1951 = ~pi014 & n333;
  assign n1952 = n1950 & n1951;
  assign n1953 = n316 & n515;
  assign n1954 = n233 & n461;
  assign n1955 = n1953 & n1954;
  assign n1956 = ~n1952 & ~n1955;
  assign n1957 = n316 & n463;
  assign n1958 = n1956 & ~n1957;
  assign n1959 = n687 & ~n1834;
  assign n1960 = n1958 & ~n1959;
  assign n1961 = ~n756 & n1960;
  assign n1962 = ~n1949 & n1961;
  assign n1963 = n1948 & n1962;
  assign n1964 = ~n1043 & ~n1307;
  assign n1965 = ~n1043 & n1302;
  assign n1966 = ~pi002 & n1551;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = ~n1964 & n1967;
  assign n1969 = n332 & n1703;
  assign n1970 = n333 & n1969;
  assign n1971 = ~n1900 & ~n1970;
  assign n1972 = ~pi011 & ~n1971;
  assign n1973 = ~pi008 & n892;
  assign n1974 = pi015 & n1973;
  assign n1975 = n1951 & n1974;
  assign n1976 = pi011 & n1975;
  assign n1977 = ~pi012 & n1185;
  assign n1978 = ~pi015 & n984;
  assign n1979 = ~n812 & ~n1978;
  assign n1980 = pi011 & ~n1979;
  assign n1981 = ~n702 & ~n1980;
  assign n1982 = ~n1977 & n1981;
  assign n1983 = n1973 & ~n1982;
  assign n1984 = ~n1976 & ~n1983;
  assign n1985 = ~n1972 & n1984;
  assign n1986 = n518 & n927;
  assign n1987 = n1089 & n1986;
  assign n1988 = ~n928 & ~n1987;
  assign n1989 = n779 & n1370;
  assign n1990 = n1988 & ~n1989;
  assign n1991 = pi014 & n865;
  assign n1992 = n1735 & n1991;
  assign n1993 = n1261 & n1992;
  assign n1994 = n1990 & ~n1993;
  assign n1995 = n1985 & n1994;
  assign n1996 = n1968 & n1995;
  assign n1997 = n1963 & n1996;
  assign n1998 = n784 & n1834;
  assign n1999 = n1262 & n1998;
  assign n2000 = ~pi043 & ~pi068;
  assign n2001 = ~pi044 & ~pi067;
  assign n2002 = n2000 & n2001;
  assign n2003 = pi042 & n2002;
  assign n2004 = n1999 & n2003;
  assign n2005 = ~pi008 & ~n458;
  assign n2006 = n979 & n2005;
  assign n2007 = n779 & n2006;
  assign n2008 = ~pi042 & n1999;
  assign n2009 = pi044 & n2000;
  assign n2010 = pi067 & n2009;
  assign n2011 = n2008 & n2010;
  assign n2012 = pi068 & n2001;
  assign n2013 = pi043 & n2012;
  assign n2014 = n2008 & n2013;
  assign n2015 = ~n2011 & ~n2014;
  assign n2016 = ~n2007 & n2015;
  assign n2017 = ~n2004 & n2016;
  assign n2018 = ~n824 & n2017;
  assign n2019 = pi005 & n1199;
  assign n2020 = n353 & n2019;
  assign n2021 = n343 & n471;
  assign n2022 = n353 & n678;
  assign n2023 = n2021 & n2022;
  assign n2024 = n1785 & n2022;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~n2020 & n2025;
  assign n2027 = n1400 & n1723;
  assign n2028 = n2026 & ~n2027;
  assign n2029 = n462 & n690;
  assign n2030 = pi014 & n691;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = n2028 & n2031;
  assign n2033 = n2018 & n2032;
  assign n2034 = n1997 & n2033;
  assign po07 = ~n1913 | ~n2034;
  assign n2036 = n583 & n934;
  assign n2037 = ~n1384 & ~n2036;
  assign n2038 = n1192 & n2037;
  assign n2039 = n495 & n592;
  assign n2040 = n335 & n2005;
  assign n2041 = ~n1719 & ~n2040;
  assign n2042 = n317 & ~n2041;
  assign n2043 = n2039 & n2042;
  assign n2044 = n1063 & ~n1936;
  assign n2045 = n1869 & n2044;
  assign n2046 = ~n1518 & ~n2045;
  assign n2047 = n676 & n1411;
  assign n2048 = n2046 & ~n2047;
  assign n2049 = ~n2043 & n2048;
  assign n2050 = n337 & n496;
  assign n2051 = pi004 & ~pi108;
  assign n2052 = n336 & n1063;
  assign n2053 = ~n2051 & n2052;
  assign n2054 = ~n2050 & ~n2053;
  assign n2055 = n284 & ~n2054;
  assign n2056 = ~n383 & n1124;
  assign n2057 = n408 & n2056;
  assign n2058 = ~n2055 & ~n2057;
  assign n2059 = n2049 & n2058;
  assign n2060 = ~n1101 & n2059;
  assign n2061 = n709 & n865;
  assign n2062 = n233 & n2061;
  assign n2063 = n458 & n2062;
  assign n2064 = ~n916 & ~n2063;
  assign n2065 = pi011 & ~n2064;
  assign n2066 = n398 & ~n2065;
  assign n2067 = n2060 & n2066;
  assign n2068 = ~pi060 & n1060;
  assign n2069 = ~pi045 & n1324;
  assign n2070 = ~pi045 & n404;
  assign n2071 = n282 & ~n2070;
  assign n2072 = ~n2069 & ~n2071;
  assign po27 = n2068 & ~n2072;
  assign n2074 = pi012 & n863;
  assign n2075 = ~n1184 & ~n2074;
  assign n2076 = n1263 & ~n2075;
  assign n2077 = ~po27 & ~n2076;
  assign n2078 = pi010 & n769;
  assign n2079 = ~n765 & ~n2078;
  assign n2080 = n702 & ~n2079;
  assign n2081 = ~n383 & n1538;
  assign n2082 = pi031 & ~pi034;
  assign n2083 = ~n693 & n2082;
  assign n2084 = ~n2081 & ~n2083;
  assign n2085 = ~n2080 & n2084;
  assign n2086 = n2077 & n2085;
  assign n2087 = n2067 & n2086;
  assign n2088 = ~pi015 & n1478;
  assign n2089 = pi008 & n510;
  assign n2090 = n416 & n2089;
  assign n2091 = n2088 & n2090;
  assign n2092 = ~pi001 & n826;
  assign n2093 = ~pi000 & n2092;
  assign n2094 = n337 & n2093;
  assign n2095 = ~pi001 & n694;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = n949 & n1285;
  assign n2098 = n2096 & ~n2097;
  assign n2099 = ~n2091 & n2098;
  assign n2100 = n357 & n2061;
  assign n2101 = ~pi014 & n2100;
  assign n2102 = n233 & n1389;
  assign n2103 = pi015 & n2102;
  assign n2104 = n274 & n460;
  assign n2105 = ~n284 & n399;
  assign n2106 = n2104 & ~n2105;
  assign n2107 = ~pi004 & n2106;
  assign n2108 = ~n2103 & ~n2107;
  assign n2109 = ~n2101 & n2108;
  assign n2110 = n982 & n1835;
  assign n2111 = ~n233 & ~n333;
  assign n2112 = n690 & ~n984;
  assign n2113 = ~n654 & n2112;
  assign n2114 = ~n2111 & n2113;
  assign n2115 = ~n2110 & ~n2114;
  assign n2116 = n284 & n848;
  assign n2117 = n1158 & n2116;
  assign n2118 = n592 & n685;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = ~n1647 & n2119;
  assign n2121 = ~n316 & ~n591;
  assign n2122 = n593 & ~n2121;
  assign n2123 = ~n946 & ~n2122;
  assign n2124 = ~n383 & ~n2123;
  assign n2125 = ~n853 & ~n2124;
  assign n2126 = n591 & n1090;
  assign n2127 = pi039 & n284;
  assign n2128 = n343 & n2039;
  assign n2129 = n2127 & n2128;
  assign n2130 = n597 & n1769;
  assign n2131 = n424 & n2130;
  assign n2132 = ~n2129 & ~n2131;
  assign n2133 = ~n2126 & n2132;
  assign n2134 = n2125 & n2133;
  assign n2135 = n2120 & n2134;
  assign n2136 = n2115 & n2135;
  assign n2137 = n2109 & n2136;
  assign n2138 = n284 & n1835;
  assign n2139 = n686 & n2138;
  assign n2140 = n688 & ~n2082;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~pi124 & ~n2141;
  assign n2143 = ~pi001 & ~pi006;
  assign n2144 = n268 & n2143;
  assign n2145 = n495 & n2144;
  assign n2146 = n2127 & n2145;
  assign n2147 = ~pi007 & n2146;
  assign n2148 = n336 & n2039;
  assign n2149 = n2127 & n2148;
  assign n2150 = ~n2147 & ~n2149;
  assign n2151 = ~n2142 & n2150;
  assign n2152 = n2137 & n2151;
  assign n2153 = n2099 & n2152;
  assign n2154 = n2087 & n2153;
  assign n2155 = n641 & n2154;
  assign n2156 = n2038 & n2155;
  assign n2157 = ~n427 & n624;
  assign n2158 = ~n649 & n2157;
  assign n2159 = n515 & n701;
  assign n2160 = n333 & n2159;
  assign n2161 = n462 & n937;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = ~pi011 & ~n2162;
  assign n2164 = ~n951 & ~n2163;
  assign n2165 = n2158 & n2164;
  assign n2166 = n568 & n2165;
  assign n2167 = n408 & n1065;
  assign n2168 = ~n1064 & ~n2167;
  assign n2169 = n354 & ~n2168;
  assign n2170 = n805 & n974;
  assign n2171 = n720 & ~n2170;
  assign n2172 = ~n2169 & n2171;
  assign n2173 = n510 & n779;
  assign n2174 = n1209 & n2173;
  assign n2175 = ~pi008 & n2174;
  assign n2176 = n233 & n1703;
  assign n2177 = n766 & n2176;
  assign n2178 = ~n2175 & ~n2177;
  assign n2179 = n274 & n494;
  assign n2180 = n423 & n2179;
  assign n2181 = ~pi006 & n2180;
  assign n2182 = ~pi002 & n2181;
  assign n2183 = n2178 & ~n2182;
  assign n2184 = n230 & n1473;
  assign n2185 = n339 & n2173;
  assign n2186 = n358 & n2185;
  assign n2187 = ~n2184 & ~n2186;
  assign n2188 = n2183 & n2187;
  assign n2189 = n2172 & n2188;
  assign n2190 = pi045 & n1060;
  assign n2191 = pi060 & n2190;
  assign n2192 = n908 & n2138;
  assign n2193 = n923 & n2192;
  assign n2194 = n370 & n1806;
  assign n2195 = pi007 & n1891;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = ~n2193 & n2196;
  assign n2198 = ~n2191 & n2197;
  assign n2199 = n432 & n1412;
  assign n2200 = n588 & n661;
  assign n2201 = n482 & n2200;
  assign n2202 = ~n2199 & ~n2201;
  assign n2203 = pi015 & n579;
  assign n2204 = n780 & n2203;
  assign n2205 = n333 & n2204;
  assign n2206 = pi015 & n1090;
  assign n2207 = n269 & n2206;
  assign n2208 = ~n2205 & ~n2207;
  assign n2209 = ~n1677 & n2208;
  assign n2210 = n2202 & n2209;
  assign n2211 = n2198 & n2210;
  assign n2212 = n2189 & n2211;
  assign n2213 = ~n381 & ~n421;
  assign n2214 = n284 & n954;
  assign n2215 = ~pi057 & n2214;
  assign n2216 = n574 & n1724;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = n2213 & n2217;
  assign n2219 = n408 & n1278;
  assign n2220 = n551 & n2219;
  assign n2221 = ~n1387 & ~n2220;
  assign n2222 = n387 & n1863;
  assign n2223 = n2221 & ~n2222;
  assign n2224 = n483 & n1667;
  assign n2225 = ~n383 & n1006;
  assign n2226 = ~pi006 & n2225;
  assign n2227 = n251 & n586;
  assign n2228 = n1126 & n2227;
  assign n2229 = n472 & n1777;
  assign n2230 = n2228 & n2229;
  assign n2231 = ~n2226 & ~n2230;
  assign n2232 = ~n1242 & n2231;
  assign n2233 = ~n2224 & n2232;
  assign n2234 = n2223 & n2233;
  assign n2235 = n776 & n805;
  assign n2236 = n777 & n2159;
  assign n2237 = n974 & n1734;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~n2235 & n2238;
  assign n2240 = n2234 & n2239;
  assign n2241 = n2218 & n2240;
  assign n2242 = n284 & ~n350;
  assign n2243 = n1153 & n1785;
  assign n2244 = n755 & n1149;
  assign n2245 = ~pi027 & n1149;
  assign n2246 = n1397 & n2245;
  assign n2247 = ~n2244 & ~n2246;
  assign n2248 = ~n2243 & n2247;
  assign n2249 = ~n2242 & n2248;
  assign n2250 = n357 & n2203;
  assign n2251 = n417 & n2250;
  assign n2252 = ~pi013 & n2251;
  assign n2253 = n315 & n791;
  assign n2254 = n2089 & n2253;
  assign n2255 = ~n689 & ~n2254;
  assign n2256 = n574 & ~n2255;
  assign n2257 = ~pi001 & n1552;
  assign n2258 = ~pi007 & n2257;
  assign n2259 = ~pi003 & n2258;
  assign n2260 = ~n2092 & ~n2259;
  assign n2261 = n346 & ~n2260;
  assign n2262 = ~pi031 & n695;
  assign n2263 = ~pi034 & n695;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = ~n2261 & n2264;
  assign n2266 = ~n2256 & n2265;
  assign n2267 = ~n2252 & n2266;
  assign n2268 = n284 & n710;
  assign n2269 = n1393 & n2268;
  assign n2270 = n384 & n730;
  assign n2271 = ~pi016 & n2270;
  assign n2272 = n482 & n2271;
  assign n2273 = ~n2269 & ~n2272;
  assign n2274 = n570 & n881;
  assign n2275 = n855 & n2271;
  assign n2276 = ~n2274 & ~n2275;
  assign n2277 = n2273 & n2276;
  assign n2278 = n577 & n2277;
  assign n2279 = n2267 & n2278;
  assign n2280 = pi100 & n1210;
  assign n2281 = n2279 & ~n2280;
  assign n2282 = n2249 & n2281;
  assign n2283 = n2241 & n2282;
  assign n2284 = n2212 & n2283;
  assign n2285 = n406 & n408;
  assign n2286 = n1619 & n2285;
  assign n2287 = ~n667 & ~n2286;
  assign n2288 = n234 & n934;
  assign n2289 = n935 & n2288;
  assign n2290 = ~pi027 & n2289;
  assign n2291 = pi014 & n905;
  assign n2292 = n547 & n2291;
  assign n2293 = pi011 & n2292;
  assign n2294 = ~n2290 & ~n2293;
  assign n2295 = n2287 & n2294;
  assign n2296 = ~n906 & ~n2291;
  assign n2297 = n926 & ~n2296;
  assign n2298 = pi007 & n1893;
  assign n2299 = ~pi012 & n815;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = n802 & ~n2300;
  assign n2302 = ~n2297 & ~n2301;
  assign n2303 = pi021 & n267;
  assign n2304 = ~n1599 & ~n2303;
  assign n2305 = pi018 & ~n2304;
  assign n2306 = ~n1360 & ~n1785;
  assign n2307 = n2305 & ~n2306;
  assign n2308 = n1728 & n2128;
  assign n2309 = ~pi119 & n2308;
  assign n2310 = ~pi110 & n269;
  assign n2311 = n1400 & n2310;
  assign n2312 = n1728 & n2311;
  assign n2313 = ~n2309 & ~n2312;
  assign n2314 = ~n955 & n2313;
  assign n2315 = n1728 & n2148;
  assign n2316 = ~pi118 & n2315;
  assign n2317 = n610 & n1625;
  assign n2318 = n533 & n1096;
  assign n2319 = n392 & n2318;
  assign n2320 = ~n2317 & ~n2319;
  assign n2321 = ~n2316 & n2320;
  assign n2322 = n2314 & n2321;
  assign n2323 = ~n2307 & n2322;
  assign n2324 = n2302 & n2323;
  assign n2325 = n2295 & n2324;
  assign n2326 = n2284 & n2325;
  assign n2327 = n2166 & n2326;
  assign po08 = ~n2156 | ~n2327;
  assign n2329 = n873 & n1224;
  assign n2330 = n508 & n700;
  assign n2331 = n926 & n2330;
  assign n2332 = n803 & n865;
  assign n2333 = ~pi009 & n2332;
  assign n2334 = pi013 & pi014;
  assign n2335 = n511 & ~n2334;
  assign n2336 = n2333 & n2335;
  assign n2337 = ~n2331 & ~n2336;
  assign n2338 = ~n2329 & n2337;
  assign n2339 = pi002 & n561;
  assign n2340 = ~n2258 & ~n2339;
  assign n2341 = pi004 & ~n2340;
  assign n2342 = ~n399 & n2341;
  assign n2343 = n2338 & ~n2342;
  assign n2344 = ~n1477 & ~n2074;
  assign n2345 = n867 & ~n2344;
  assign n2346 = n1998 & n2333;
  assign n2347 = pi015 & n2346;
  assign n2348 = ~n1612 & ~n2347;
  assign n2349 = ~n2345 & n2348;
  assign n2350 = n2343 & n2349;
  assign n2351 = n543 & n1607;
  assign n2352 = pi013 & n866;
  assign n2353 = n789 & n2352;
  assign n2354 = pi010 & n2353;
  assign n2355 = ~n2351 & ~n2354;
  assign n2356 = ~pi123 & ~n2355;
  assign n2357 = ~n1301 & ~n1549;
  assign n2358 = pi002 & n574;
  assign n2359 = n2179 & n2358;
  assign n2360 = n224 & n2359;
  assign n2361 = n2357 & ~n2360;
  assign n2362 = pi002 & n2180;
  assign n2363 = n2361 & ~n2362;
  assign n2364 = ~n2356 & n2363;
  assign n2365 = n2350 & n2364;
  assign n2366 = n388 & n843;
  assign n2367 = ~n841 & ~n2366;
  assign n2368 = pi022 & ~n2367;
  assign n2369 = ~pi015 & n2298;
  assign n2370 = n1889 & n2369;
  assign n2371 = ~pi003 & pi007;
  assign n2372 = n2257 & n2371;
  assign n2373 = n1547 & n2372;
  assign n2374 = pi002 & n1847;
  assign n2375 = n337 & n2374;
  assign n2376 = ~n2373 & ~n2375;
  assign n2377 = ~n2370 & n2376;
  assign n2378 = n866 & n1876;
  assign n2379 = n803 & n1977;
  assign n2380 = n708 & n1184;
  assign n2381 = n547 & n1225;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = ~n2379 & n2382;
  assign n2384 = n1991 & ~n2383;
  assign n2385 = ~n2378 & ~n2384;
  assign n2386 = n2377 & n2385;
  assign n2387 = ~n2368 & n2386;
  assign n2388 = n480 & n1525;
  assign n2389 = n411 & n843;
  assign n2390 = n843 & n1600;
  assign n2391 = ~pi020 & n2390;
  assign n2392 = n1846 & n2358;
  assign n2393 = n345 & n1552;
  assign n2394 = ~n2392 & ~n2393;
  assign n2395 = n592 & ~n2394;
  assign n2396 = ~n2391 & ~n2395;
  assign n2397 = ~n2389 & n2396;
  assign n2398 = ~n2388 & n2397;
  assign n2399 = n2387 & n2398;
  assign n2400 = n809 & n865;
  assign n2401 = n744 & ~n2400;
  assign n2402 = pi011 & n1226;
  assign n2403 = n804 & n1224;
  assign n2404 = ~n462 & ~n800;
  assign n2405 = n2403 & ~n2404;
  assign n2406 = ~n2402 & ~n2405;
  assign n2407 = n274 & n2392;
  assign n2408 = ~pi122 & n2407;
  assign n2409 = n336 & n2259;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n388 & ~n644;
  assign n2412 = ~n383 & n836;
  assign n2413 = ~n2411 & n2412;
  assign n2414 = n2410 & ~n2413;
  assign n2415 = n2406 & n2414;
  assign n2416 = n2401 & n2415;
  assign n2417 = n2399 & n2416;
  assign po09 = ~n2365 | ~n2417;
  assign n2419 = n619 & n1312;
  assign n2420 = ~n1344 & ~n2419;
  assign n2421 = n619 & n999;
  assign n2422 = ~n1003 & n2421;
  assign n2423 = n619 & n961;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = n2420 & n2424;
  assign n2426 = n511 & n871;
  assign n2427 = n354 & n2426;
  assign n2428 = n779 & n2427;
  assign n2429 = ~n915 & n2428;
  assign n2430 = ~n939 & ~n2429;
  assign n2431 = n512 & n937;
  assign n2432 = n2430 & ~n2431;
  assign n2433 = n804 & n974;
  assign n2434 = ~n2298 & ~n2433;
  assign n2435 = n234 & ~n2434;
  assign n2436 = ~n818 & ~n2435;
  assign n2437 = n811 & ~n2436;
  assign n2438 = pi027 & n2437;
  assign n2439 = pi015 & n936;
  assign n2440 = n702 & n2439;
  assign n2441 = ~n2438 & ~n2440;
  assign n2442 = n2432 & n2441;
  assign n2443 = n2425 & n2442;
  assign n2444 = n234 & n801;
  assign n2445 = n978 & n2444;
  assign n2446 = n708 & n2445;
  assign n2447 = n717 & n969;
  assign n2448 = n949 & n965;
  assign n2449 = ~pi037 & n2448;
  assign n2450 = n1346 & n2449;
  assign n2451 = ~n2447 & ~n2450;
  assign n2452 = n354 & n973;
  assign n2453 = pi035 & n970;
  assign n2454 = n1869 & n2453;
  assign n2455 = ~n2452 & ~n2454;
  assign n2456 = n2451 & n2455;
  assign n2457 = ~n2446 & n2456;
  assign n2458 = n354 & n632;
  assign n2459 = n729 & n2458;
  assign n2460 = n2457 & ~n2459;
  assign n2461 = n516 & n978;
  assign n2462 = n710 & n2461;
  assign n2463 = ~pi013 & n924;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = n1991 & n2369;
  assign n2466 = n918 & ~n2465;
  assign n2467 = n2464 & n2466;
  assign n2468 = n905 & n1186;
  assign n2469 = pi011 & n701;
  assign n2470 = ~n712 & ~n2469;
  assign n2471 = ~n2468 & n2470;
  assign n2472 = n1237 & n2471;
  assign n2473 = n2467 & n2472;
  assign n2474 = pi012 & n2444;
  assign n2475 = ~n817 & n2474;
  assign n2476 = n462 & n804;
  assign n2477 = n2444 & n2476;
  assign n2478 = ~n2475 & ~n2477;
  assign n2479 = n776 & n2334;
  assign n2480 = n709 & n2479;
  assign n2481 = ~n2298 & ~n2480;
  assign n2482 = n914 & ~n2481;
  assign n2483 = n707 & n2482;
  assign n2484 = n2478 & ~n2483;
  assign n2485 = n333 & n922;
  assign n2486 = pi007 & n2485;
  assign n2487 = n1889 & n2486;
  assign n2488 = pi009 & n2487;
  assign n2489 = ~pi015 & n2488;
  assign n2490 = n337 & n2372;
  assign n2491 = n777 & n2061;
  assign n2492 = n230 & n2257;
  assign po48 = ~n2371 & n2492;
  assign n2494 = ~n2491 & ~po48;
  assign n2495 = ~n2490 & n2494;
  assign n2496 = ~n2489 & n2495;
  assign n2497 = n2484 & n2496;
  assign n2498 = n235 & n905;
  assign n2499 = ~pi011 & n2498;
  assign n2500 = n368 & n1452;
  assign n2501 = n471 & n1383;
  assign n2502 = n269 & n2501;
  assign n2503 = ~n2500 & ~n2502;
  assign n2504 = ~n1345 & n2503;
  assign n2505 = ~n2499 & n2504;
  assign n2506 = pi123 & ~n2355;
  assign n2507 = n2505 & ~n2506;
  assign n2508 = n2497 & n2507;
  assign n2509 = n2473 & n2508;
  assign n2510 = n2460 & n2509;
  assign po10 = ~n2443 | ~n2510;
  assign n2512 = n734 & n2229;
  assign n2513 = n230 & n471;
  assign n2514 = n433 & n2513;
  assign n2515 = ~n2271 & ~n2514;
  assign n2516 = n553 & ~n2515;
  assign n2517 = n230 & n469;
  assign n2518 = n1562 & n2517;
  assign n2519 = n949 & n2517;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = ~n1196 & n2520;
  assign n2522 = ~n2516 & n2521;
  assign n2523 = ~n857 & n2522;
  assign n2524 = ~n2512 & n2523;
  assign n2525 = ~pi013 & n867;
  assign n2526 = ~n789 & n2525;
  assign n2527 = ~n1153 & ~n1201;
  assign n2528 = n735 & ~n2527;
  assign n2529 = ~n2526 & ~n2528;
  assign n2530 = n1594 & n2412;
  assign n2531 = ~n1632 & ~n2374;
  assign n2532 = ~pi007 & ~n2531;
  assign n2533 = n346 & n2532;
  assign n2534 = n316 & n2257;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = ~n2530 & n2535;
  assign n2537 = n408 & n1451;
  assign n2538 = n374 & n732;
  assign n2539 = pi019 & n2538;
  assign n2540 = ~n2537 & ~n2539;
  assign n2541 = n2536 & n2540;
  assign n2542 = n1331 & n1414;
  assign n2543 = ~n870 & ~n2542;
  assign n2544 = ~pi022 & n841;
  assign n2545 = n725 & n752;
  assign n2546 = ~pi022 & n2545;
  assign n2547 = ~n2544 & ~n2546;
  assign n2548 = n533 & n1359;
  assign n2549 = n373 & n2548;
  assign n2550 = ~n775 & ~n2549;
  assign n2551 = n729 & n2271;
  assign n2552 = n2550 & ~n2551;
  assign n2553 = n2547 & n2552;
  assign n2554 = n2543 & n2553;
  assign n2555 = n2541 & n2554;
  assign n2556 = n2529 & n2555;
  assign n2557 = n2524 & n2556;
  assign n2558 = n374 & n2514;
  assign n2559 = ~pi022 & n1610;
  assign n2560 = n230 & n2559;
  assign n2561 = n369 & n2560;
  assign n2562 = ~n2558 & ~n2561;
  assign n2563 = pi021 & ~n2562;
  assign n2564 = n469 & n723;
  assign n2565 = n1278 & n2513;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = n678 & n2271;
  assign n2568 = n678 & n1126;
  assign n2569 = n394 & n2568;
  assign n2570 = ~n2567 & ~n2569;
  assign n2571 = n2566 & n2570;
  assign n2572 = n384 & n1610;
  assign n2573 = n394 & n1599;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n469 & ~n2574;
  assign n2576 = n1414 & n2513;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = n2571 & n2577;
  assign n2579 = n1108 & n1359;
  assign n2580 = n230 & n2579;
  assign n2581 = ~pi017 & n2580;
  assign n2582 = n2578 & ~n2581;
  assign n2583 = ~n2563 & n2582;
  assign n2584 = pi016 & n856;
  assign n2585 = n375 & n2584;
  assign n2586 = ~n1198 & ~n2585;
  assign n2587 = n725 & n1599;
  assign n2588 = n2586 & ~n2587;
  assign n2589 = ~pi082 & n952;
  assign n2590 = n2588 & ~n2589;
  assign n2591 = ~n1610 & ~n2303;
  assign n2592 = pi020 & ~n2591;
  assign n2593 = ~n774 & ~n2592;
  assign n2594 = ~n958 & n2593;
  assign n2595 = n394 & ~n2594;
  assign n2596 = n394 & n1201;
  assign n2597 = n230 & n569;
  assign n2598 = ~n2596 & ~n2597;
  assign n2599 = ~pi020 & ~n2598;
  assign n2600 = ~n2595 & ~n2599;
  assign n2601 = n661 & ~n2600;
  assign n2602 = n277 & n409;
  assign n2603 = n472 & n1408;
  assign n2604 = ~n678 & ~n958;
  assign n2605 = ~n2603 & n2604;
  assign n2606 = n661 & ~n2605;
  assign n2607 = ~n2602 & ~n2606;
  assign n2608 = n384 & ~n2607;
  assign n2609 = n966 & n2513;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = ~n2601 & n2610;
  assign n2612 = n709 & n1992;
  assign n2613 = n2611 & ~n2612;
  assign n2614 = ~n662 & ~n1778;
  assign n2615 = n386 & ~n2614;
  assign n2616 = n2613 & ~n2615;
  assign n2617 = n2590 & n2616;
  assign n2618 = n2583 & n2617;
  assign po11 = ~n2557 | ~n2618;
  assign n2620 = n274 & n1552;
  assign n2621 = n408 & n1741;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = n480 & ~n2622;
  assign n2624 = n509 & n1893;
  assign n2625 = n728 & ~n2624;
  assign n2626 = ~n2623 & n2625;
  assign n2627 = n333 & n814;
  assign n2628 = n1889 & n2627;
  assign n2629 = n334 & n766;
  assign n2630 = n517 & n2629;
  assign n2631 = ~n2488 & ~n2630;
  assign n2632 = ~n2628 & n2631;
  assign n2633 = pi015 & ~n2632;
  assign n2634 = n812 & n2352;
  assign n2635 = pi011 & n2634;
  assign n2636 = ~pi022 & n2366;
  assign n2637 = n1552 & n2144;
  assign n2638 = n1020 & n1889;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = pi007 & ~n2639;
  assign n2641 = ~n2636 & ~n2640;
  assign n2642 = ~n2635 & n2641;
  assign n2643 = ~n2633 & n2642;
  assign po12 = ~n2626 | ~n2643;
  assign n2645 = pi124 & ~n2141;
  assign n2646 = n1785 & n2305;
  assign n2647 = n692 & ~n2082;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = ~n2645 & n2648;
  assign n2650 = n690 & n2138;
  assign n2651 = ~n2118 & ~n2650;
  assign n2652 = ~n2244 & n2651;
  assign n2653 = pi064 & n2047;
  assign n2654 = ~pi017 & n2653;
  assign n2655 = ~n2030 & ~n2654;
  assign n2656 = n2652 & n2655;
  assign po13 = ~n2649 | ~n2656;
  assign n2658 = ~pi011 & ~n1988;
  assign n2659 = ~n456 & n1761;
  assign n2660 = ~pi019 & ~n2659;
  assign n2661 = ~n1905 & n2025;
  assign n2662 = n570 & n1562;
  assign n2663 = pi023 & n1879;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = n2661 & n2664;
  assign n2666 = ~n2660 & n2665;
  assign n2667 = ~n2658 & n2666;
  assign n2668 = n234 & n1838;
  assign n2669 = pi008 & n2668;
  assign n2670 = ~n1807 & ~n2669;
  assign n2671 = ~n1363 & n2670;
  assign n2672 = ~n716 & n1372;
  assign n2673 = n224 & n1875;
  assign n2674 = n982 & n2673;
  assign n2675 = ~n2672 & ~n2674;
  assign n2676 = n1985 & n2675;
  assign n2677 = n2671 & n2676;
  assign n2678 = n1290 & n2288;
  assign n2679 = ~n1529 & ~n2678;
  assign n2680 = n589 & n752;
  assign n2681 = ~n1648 & ~n2680;
  assign n2682 = n444 & n773;
  assign n2683 = n2681 & ~n2682;
  assign n2684 = n1696 & n2683;
  assign n2685 = ~n687 & ~n1091;
  assign n2686 = ~pi015 & ~n2685;
  assign n2687 = n317 & n2206;
  assign n2688 = ~pi011 & n1749;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2686 & n2689;
  assign n2691 = pi014 & ~n2690;
  assign n2692 = n2684 & ~n2691;
  assign n2693 = n2679 & n2692;
  assign n2694 = ~n1070 & n1705;
  assign n2695 = ~pi019 & n2694;
  assign n2696 = n284 & n2019;
  assign n2697 = pi004 & n2696;
  assign n2698 = ~pi006 & n1955;
  assign n2699 = ~n2225 & ~n2698;
  assign n2700 = ~n2697 & n2699;
  assign n2701 = n1166 & n1176;
  assign n2702 = ~n1318 & ~n2319;
  assign n2703 = ~n2701 & n2702;
  assign n2704 = n2700 & n2703;
  assign n2705 = ~n2695 & n2704;
  assign n2706 = n511 & n1183;
  assign n2707 = ~n511 & n1734;
  assign n2708 = ~n2706 & ~n2707;
  assign n2709 = ~pi013 & ~n2708;
  assign n2710 = n432 & n840;
  assign n2711 = ~n385 & n2710;
  assign n2712 = ~n2709 & ~n2711;
  assign n2713 = n1711 & n2712;
  assign n2714 = n2705 & n2713;
  assign n2715 = n2693 & n2714;
  assign n2716 = n2677 & n2715;
  assign n2717 = ~n1935 & n1939;
  assign n2718 = n616 & n1166;
  assign n2719 = ~pi113 & n1169;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = ~n2717 & n2720;
  assign n2722 = n704 & n779;
  assign n2723 = n2426 & n2722;
  assign n2724 = n758 & n1561;
  assign n2725 = n372 & n2724;
  assign n2726 = ~n2723 & ~n2725;
  assign n2727 = ~n1264 & n2726;
  assign n2728 = n1288 & n2727;
  assign n2729 = ~pi004 & ~pi006;
  assign n2730 = n1840 & n2729;
  assign n2731 = ~n1712 & ~n2730;
  assign n2732 = n2728 & n2731;
  assign n2733 = ~pi011 & n1903;
  assign n2734 = ~n1532 & ~n2733;
  assign n2735 = ~pi021 & n1384;
  assign n2736 = n747 & n754;
  assign n2737 = ~n1546 & ~n2736;
  assign n2738 = ~n2735 & n2737;
  assign n2739 = n2734 & n2738;
  assign n2740 = n2732 & n2739;
  assign n2741 = n2721 & n2740;
  assign n2742 = n376 & n484;
  assign n2743 = ~n664 & ~n2742;
  assign n2744 = n432 & ~n2743;
  assign n2745 = ~pi022 & n2224;
  assign n2746 = n333 & n515;
  assign n2747 = n690 & n2746;
  assign n2748 = n1874 & ~n2747;
  assign n2749 = ~n2745 & n2748;
  assign n2750 = ~n2744 & n2749;
  assign n2751 = n626 & n758;
  assign n2752 = n647 & n1835;
  assign n2753 = ~n1652 & ~n2752;
  assign n2754 = ~n2751 & n2753;
  assign n2755 = n2750 & n2754;
  assign n2756 = n2164 & n2755;
  assign n2757 = n2741 & n2756;
  assign n2758 = n2716 & n2757;
  assign n2759 = n2667 & n2758;
  assign n2760 = ~n1856 & n2221;
  assign n2761 = n1898 & n2760;
  assign n2762 = ~pi027 & n1398;
  assign n2763 = n892 & n1209;
  assign n2764 = n1410 & n1459;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = ~n1755 & n2765;
  assign n2767 = ~n2762 & n2766;
  assign n2768 = ~n383 & n1050;
  assign n2769 = ~n1222 & ~n2768;
  assign n2770 = n2767 & n2769;
  assign n2771 = n2761 & n2770;
  assign n2772 = ~n625 & ~n627;
  assign n2773 = n343 & ~n2772;
  assign n2774 = ~n1107 & ~n2773;
  assign n2775 = ~n981 & n2774;
  assign n2776 = ~n1070 & ~n2775;
  assign n2777 = n726 & n1303;
  assign n2778 = ~n1043 & n2777;
  assign n2779 = n1414 & n1864;
  assign n2780 = n443 & n470;
  assign n2781 = pi019 & n2780;
  assign n2782 = n1241 & ~n1655;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = ~n2779 & n2783;
  assign n2785 = pi015 & n1476;
  assign n2786 = ~n2199 & ~n2785;
  assign n2787 = n2784 & n2786;
  assign n2788 = ~n2778 & n2787;
  assign n2789 = ~n2776 & n2788;
  assign n2790 = pi122 & ~n1937;
  assign n2791 = ~n1747 & ~n2790;
  assign n2792 = n1934 & n2791;
  assign n2793 = ~n1213 & n1330;
  assign n2794 = n1789 & n2793;
  assign n2795 = n2792 & n2794;
  assign n2796 = ~n1174 & n1439;
  assign n2797 = n780 & n1478;
  assign n2798 = n978 & n2722;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = ~pi010 & ~n2799;
  assign n2801 = n473 & n661;
  assign n2802 = ~n844 & ~n2801;
  assign n2803 = n588 & ~n2802;
  assign n2804 = ~n2800 & ~n2803;
  assign n2805 = ~n915 & n1259;
  assign n2806 = ~n458 & n2805;
  assign n2807 = ~n1636 & ~n2806;
  assign n2808 = n2804 & n2807;
  assign n2809 = n2796 & n2808;
  assign n2810 = n230 & n1840;
  assign n2811 = n1450 & ~n2810;
  assign n2812 = ~pi089 & n2668;
  assign n2813 = n2811 & ~n2812;
  assign n2814 = n1876 & n1973;
  assign n2815 = ~pi020 & ~pi021;
  assign n2816 = n1757 & ~n2815;
  assign n2817 = ~n2814 & ~n2816;
  assign n2818 = pi015 & ~n2031;
  assign n2819 = n229 & n1473;
  assign n2820 = ~n1957 & ~n2819;
  assign n2821 = ~pi015 & ~n2820;
  assign n2822 = pi014 & ~n333;
  assign n2823 = n1949 & ~n2822;
  assign n2824 = ~n1623 & ~n2823;
  assign n2825 = ~n2821 & n2824;
  assign n2826 = n1795 & n2825;
  assign n2827 = ~n2818 & n2826;
  assign n2828 = n2817 & n2827;
  assign n2829 = n2813 & n2828;
  assign n2830 = n2809 & n2829;
  assign n2831 = n2018 & n2830;
  assign n2832 = n2795 & n2831;
  assign n2833 = n2789 & n2832;
  assign n2834 = n2771 & n2833;
  assign po14 = ~n2759 | ~n2834;
  assign n2836 = n1368 & n2320;
  assign n2837 = n2794 & n2836;
  assign n2838 = ~pi007 & n1848;
  assign n2839 = n229 & n2838;
  assign n2840 = pi014 & n1949;
  assign n2841 = ~n1089 & n2729;
  assign n2842 = n1090 & n2841;
  assign n2843 = ~n2840 & ~n2842;
  assign n2844 = ~n2839 & n2843;
  assign n2845 = n705 & n1834;
  assign n2846 = ~n1735 & ~n2845;
  assign n2847 = n701 & ~n2846;
  assign n2848 = n2844 & ~n2847;
  assign n2849 = pi020 & pi021;
  assign n2850 = n375 & n2849;
  assign n2851 = ~n385 & ~n1610;
  assign n2852 = n2815 & ~n2851;
  assign n2853 = ~n2850 & ~n2852;
  assign n2854 = n734 & ~n2853;
  assign n2855 = ~pi015 & n2184;
  assign n2856 = ~n1831 & ~n2855;
  assign n2857 = ~n2854 & n2856;
  assign n2858 = n2848 & n2857;
  assign n2859 = ~n873 & ~n1225;
  assign n2860 = n1991 & ~n2859;
  assign n2861 = ~pi002 & ~n308;
  assign n2862 = ~pi005 & ~pi007;
  assign n2863 = n1085 & ~n2862;
  assign n2864 = ~n2861 & n2863;
  assign n2865 = ~n459 & n494;
  assign n2866 = ~pi001 & n2865;
  assign n2867 = ~n2864 & n2866;
  assign n2868 = ~n399 & n2861;
  assign n2869 = ~pi004 & n2868;
  assign n2870 = n2867 & ~n2869;
  assign n2871 = ~n250 & n548;
  assign n2872 = n461 & n2871;
  assign n2873 = ~n2121 & n2872;
  assign n2874 = ~n2870 & ~n2873;
  assign n2875 = n1956 & n2874;
  assign n2876 = ~n894 & n2875;
  assign n2877 = ~n2860 & n2876;
  assign n2878 = n2858 & n2877;
  assign n2879 = ~n1448 & ~n1480;
  assign n2880 = n1757 & ~n2849;
  assign n2881 = n2879 & ~n2880;
  assign n2882 = n777 & n923;
  assign n2883 = ~n2269 & ~n2882;
  assign n2884 = n2881 & n2883;
  assign n2885 = n2878 & n2884;
  assign n2886 = n701 & n934;
  assign n2887 = n1089 & n2886;
  assign n2888 = n2632 & ~n2887;
  assign n2889 = ~pi012 & n867;
  assign n2890 = ~n1442 & ~n2889;
  assign n2891 = n2888 & n2890;
  assign n2892 = n2885 & n2891;
  assign n2893 = ~n627 & ~n706;
  assign n2894 = n1426 & ~n2893;
  assign n2895 = ~n724 & ~n2615;
  assign n2896 = ~n733 & n2895;
  assign n2897 = n958 & n2271;
  assign n2898 = ~n2539 & ~n2897;
  assign n2899 = n2896 & n2898;
  assign n2900 = ~n2894 & n2899;
  assign n2901 = n2892 & n2900;
  assign n2902 = n490 & n836;
  assign n2903 = n1599 & n2902;
  assign n2904 = n2348 & ~n2903;
  assign n2905 = n1273 & n1296;
  assign n2906 = n2904 & n2905;
  assign n2907 = n2771 & n2906;
  assign n2908 = n2901 & n2907;
  assign n2909 = ~pi017 & n1695;
  assign n2910 = n462 & n927;
  assign n2911 = pi015 & n1790;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = ~n2909 & n2912;
  assign n2914 = n562 & n574;
  assign n2915 = ~n2130 & ~n2914;
  assign n2916 = ~n1095 & n2915;
  assign n2917 = n317 & n463;
  assign n2918 = n591 & n1474;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = pi015 & ~n2919;
  assign n2921 = n2100 & ~n2334;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = n2916 & n2922;
  assign n2924 = n2913 & n2923;
  assign n2925 = ~n1047 & ~po67;
  assign n2926 = ~n374 & ~n467;
  assign n2927 = n444 & ~n2926;
  assign n2928 = n2562 & ~n2927;
  assign n2929 = n2925 & n2928;
  assign n2930 = n2924 & n2929;
  assign n2931 = n354 & n633;
  assign n2932 = ~n1345 & ~n2931;
  assign n2933 = n714 & n1906;
  assign n2934 = n2932 & n2933;
  assign n2935 = n2523 & n2934;
  assign n2936 = n2930 & n2935;
  assign n2937 = n1559 & n2936;
  assign n2938 = n2033 & n2937;
  assign n2939 = n2908 & n2938;
  assign n2940 = n2837 & n2939;
  assign n2941 = ~n1259 & ~n1902;
  assign n2942 = n458 & ~n2941;
  assign n2943 = n224 & ~n1566;
  assign n2944 = ~n446 & n1640;
  assign n2945 = ~n1589 & ~n2944;
  assign n2946 = ~n2943 & n2945;
  assign n2947 = ~n2942 & n2946;
  assign n2948 = n923 & n2479;
  assign n2949 = n334 & n704;
  assign n2950 = ~n1998 & ~n2949;
  assign n2951 = pi015 & n2268;
  assign n2952 = ~n2950 & n2951;
  assign n2953 = ~n2948 & ~n2952;
  assign n2954 = n2338 & n2953;
  assign n2955 = ~n2353 & ~n2634;
  assign n2956 = pi010 & ~n2955;
  assign n2957 = n1876 & n2332;
  assign n2958 = n789 & n914;
  assign n2959 = n711 & n2958;
  assign n2960 = n1889 & n1893;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = ~n2957 & n2961;
  assign n2963 = ~n2956 & n2962;
  assign n2964 = n2954 & n2963;
  assign n2965 = ~n742 & n2611;
  assign n2966 = ~n2545 & n2550;
  assign n2967 = ~n2580 & n2966;
  assign n2968 = n2965 & n2967;
  assign n2969 = n2964 & n2968;
  assign n2970 = n2947 & n2969;
  assign n2971 = n443 & n1526;
  assign n2972 = ~n458 & n1090;
  assign n2973 = ~n2093 & ~n2972;
  assign n2974 = n230 & ~n2973;
  assign n2975 = n251 & n463;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = ~n1697 & n2976;
  assign n2978 = ~n1694 & ~n2637;
  assign n2979 = n2977 & n2978;
  assign n2980 = ~n2971 & n2979;
  assign n2981 = n953 & n2980;
  assign n2982 = n451 & ~n2586;
  assign n2983 = n1762 & n2425;
  assign n2984 = ~n2982 & n2983;
  assign n2985 = n2981 & n2984;
  assign n2986 = n2970 & n2985;
  assign n2987 = n1948 & n2986;
  assign n2988 = n2940 & n2987;
  assign n2989 = pi005 & n1575;
  assign n2990 = ~n1115 & ~n1310;
  assign n2991 = ~n2989 & n2990;
  assign n2992 = n1756 & n2021;
  assign n2993 = n482 & n1276;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = n224 & ~n2994;
  assign n2996 = n224 & n343;
  assign n2997 = n1561 & n2996;
  assign n2998 = ~pi122 & n250;
  assign n2999 = ~n1585 & ~n2998;
  assign n3000 = ~n2997 & n2999;
  assign n3001 = ~n1561 & ~n1756;
  assign n3002 = n471 & ~n3001;
  assign n3003 = ~n3000 & n3002;
  assign n3004 = ~n2995 & ~n3003;
  assign n3005 = n1778 & n1862;
  assign n3006 = ~n486 & ~n1653;
  assign n3007 = ~n3005 & n3006;
  assign n3008 = n3004 & n3007;
  assign n3009 = n392 & n2412;
  assign n3010 = n729 & n3009;
  assign n3011 = n446 & n1607;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n2391 & n3012;
  assign n3014 = pi018 & ~n3013;
  assign n3015 = n3008 & ~n3014;
  assign n3016 = n354 & n586;
  assign n3017 = pi065 & n3016;
  assign n3018 = n1070 & ~n3017;
  assign n3019 = n960 & ~n3018;
  assign n3020 = ~n1332 & ~n3019;
  assign n3021 = n224 & n1417;
  assign n3022 = ~n1636 & ~n3021;
  assign n3023 = ~n1661 & n3022;
  assign n3024 = n3020 & n3023;
  assign n3025 = n274 & n1846;
  assign n3026 = ~pi002 & ~n342;
  assign n3027 = ~n383 & ~n3026;
  assign n3028 = n3025 & n3027;
  assign n3029 = ~n1116 & n3028;
  assign n3030 = ~pi007 & n1631;
  assign n3031 = n423 & n3030;
  assign n3032 = ~n2224 & ~n3031;
  assign n3033 = ~n3029 & n3032;
  assign n3034 = n3024 & n3033;
  assign n3035 = n3015 & n3034;
  assign n3036 = n2991 & n3035;
  assign n3037 = ~n1437 & ~n1797;
  assign n3038 = ~n1071 & ~n1471;
  assign n3039 = n1319 & n3038;
  assign n3040 = n3037 & n3039;
  assign n3041 = ~n987 & ~n1070;
  assign n3042 = n1628 & ~n3041;
  assign n3043 = ~n702 & ~n1184;
  assign n3044 = n1183 & ~n3043;
  assign n3045 = ~n598 & ~n3044;
  assign n3046 = ~n2780 & n3045;
  assign n3047 = n1179 & n3046;
  assign n3048 = n3042 & n3047;
  assign n3049 = n3040 & n3048;
  assign n3050 = n1143 & ~n1767;
  assign n3051 = n455 & n3050;
  assign n3052 = n1008 & n1139;
  assign n3053 = n3051 & n3052;
  assign n3054 = ~n383 & ~n3053;
  assign n3055 = n846 & ~n1099;
  assign n3056 = ~n1597 & n3055;
  assign n3057 = ~n1079 & ~n1868;
  assign n3058 = n3056 & n3057;
  assign n3059 = n834 & n2227;
  assign n3060 = n423 & n1299;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = n1714 & n2754;
  assign n3063 = n3061 & n3062;
  assign n3064 = n3058 & n3063;
  assign n3065 = ~n3054 & n3064;
  assign n3066 = n3049 & n3065;
  assign n3067 = n3036 & n3066;
  assign n3068 = n354 & ~n1067;
  assign n3069 = ~n1706 & ~n3068;
  assign n3070 = ~n829 & n2457;
  assign n3071 = n3069 & n3070;
  assign n3072 = n1304 & n2271;
  assign n3073 = ~n385 & n387;
  assign n3074 = n735 & n3073;
  assign n3075 = ~n3072 & ~n3074;
  assign n3076 = ~n955 & n3075;
  assign n3077 = n2578 & n3076;
  assign n3078 = n2217 & n3077;
  assign n3079 = ~n1747 & n3078;
  assign n3080 = n1069 & ~n1547;
  assign n3081 = n1334 & n3080;
  assign n3082 = n638 & n1069;
  assign n3083 = ~pi061 & n3082;
  assign n3084 = ~n3081 & ~n3083;
  assign n3085 = ~n1476 & n3084;
  assign n3086 = n1252 & n3085;
  assign n3087 = n496 & n2127;
  assign n3088 = n1547 & n3087;
  assign n3089 = ~n1730 & ~n3088;
  assign n3090 = n251 & n2838;
  assign n3091 = ~pi088 & n3090;
  assign n3092 = n270 & ~n385;
  assign n3093 = n1396 & n3092;
  assign n3094 = ~n3091 & ~n3093;
  assign n3095 = ~n1482 & n3094;
  assign n3096 = n3089 & n3095;
  assign n3097 = ~n1872 & n3096;
  assign n3098 = n3086 & n3097;
  assign n3099 = n3079 & n3098;
  assign n3100 = pi015 & n1371;
  assign n3101 = ~n1720 & ~n1817;
  assign n3102 = ~n3100 & n3101;
  assign n3103 = n2675 & n3102;
  assign n3104 = n3099 & n3103;
  assign n3105 = ~n1233 & n3104;
  assign n3106 = n3071 & n3105;
  assign n3107 = n2430 & ~n2475;
  assign n3108 = n1875 & n2469;
  assign n3109 = ~pi013 & n906;
  assign n3110 = ~pi014 & n511;
  assign n3111 = n3109 & ~n3110;
  assign n3112 = ~n3108 & ~n3111;
  assign n3113 = ~n1186 & n2627;
  assign n3114 = n702 & n813;
  assign n3115 = ~n2433 & ~n3114;
  assign n3116 = ~n2299 & n3115;
  assign n3117 = ~n3113 & n3116;
  assign n3118 = n1224 & ~n3117;
  assign n3119 = n3112 & ~n3118;
  assign n3120 = n3107 & n3119;
  assign n3121 = n361 & n913;
  assign n3122 = ~n516 & ~n2958;
  assign n3123 = pi011 & ~n3122;
  assign n3124 = n913 & n3123;
  assign n3125 = ~n1704 & ~n3124;
  assign n3126 = ~n3121 & n3125;
  assign n3127 = ~n917 & n3126;
  assign n3128 = ~n2498 & n3127;
  assign n3129 = ~n2292 & n3128;
  assign n3130 = ~n2289 & n3129;
  assign n3131 = ~n816 & ~n2298;
  assign n3132 = n1224 & ~n3131;
  assign n3133 = n3130 & ~n3132;
  assign n3134 = n515 & n935;
  assign n3135 = n803 & n2444;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = n702 & ~n3136;
  assign n3138 = ~n2437 & ~n3137;
  assign n3139 = n3133 & n3138;
  assign n3140 = n3120 & n3139;
  assign n3141 = ~n1793 & ~n1901;
  assign n3142 = n1995 & n3141;
  assign n3143 = ~n2111 & n2159;
  assign n3144 = n3142 & ~n3143;
  assign n3145 = ~n2251 & n3144;
  assign n3146 = ~n897 & ~n2669;
  assign n3147 = ~n2812 & n3146;
  assign n3148 = ~n1891 & ~n2161;
  assign n3149 = n3147 & n3148;
  assign n3150 = n705 & n1718;
  assign n3151 = n700 & n3150;
  assign n3152 = n234 & n705;
  assign n3153 = n701 & n3152;
  assign n3154 = ~n3151 & ~n3153;
  assign n3155 = ~n1737 & n3154;
  assign n3156 = n3149 & n3155;
  assign n3157 = n3145 & n3156;
  assign n3158 = n3140 & n3157;
  assign n3159 = n3106 & n3158;
  assign n3160 = n3067 & n3159;
  assign po15 = ~n2988 | ~n3160;
  assign n3162 = n354 & n651;
  assign n3163 = ~n1845 & ~n3162;
  assign n3164 = n2018 & n3163;
  assign n3165 = n569 & ~n2306;
  assign n3166 = ~n422 & ~n3165;
  assign n3167 = n3164 & n3166;
  assign n3168 = ~n2286 & n3167;
  assign n3169 = ~n364 & ~n1022;
  assign n3170 = ~n1014 & n3169;
  assign n3171 = ~n257 & ~n263;
  assign n3172 = n3170 & ~n3171;
  assign n3173 = pi044 & ~pi055;
  assign n3174 = n1930 & ~n3173;
  assign n3175 = ~n1164 & n3174;
  assign n3176 = pi044 & n1930;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3172 & ~n3177;
  assign n3179 = ~pi056 & n337;
  assign n3180 = ~n528 & ~n3179;
  assign n3181 = n297 & ~n3180;
  assign n3182 = n257 & ~n1017;
  assign n3183 = ~pi122 & ~n3182;
  assign n3184 = ~n294 & ~n325;
  assign n3185 = ~n280 & n3184;
  assign n3186 = ~n3183 & n3185;
  assign n3187 = ~pi045 & ~n3186;
  assign n3188 = ~n3181 & ~n3187;
  assign n3189 = ~n3178 & n3188;
  assign n3190 = ~n1914 & ~n3175;
  assign n3191 = ~n3176 & n3190;
  assign n3192 = n1029 & ~n3191;
  assign n3193 = ~pi045 & n1074;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = n3189 & n3194;
  assign n3196 = ~pi020 & n393;
  assign n3197 = n1135 & n3196;
  assign n3198 = ~pi045 & n3197;
  assign n3199 = ~pi005 & n3198;
  assign n3200 = ~n287 & ~po27;
  assign n3201 = ~n3199 & n3200;
  assign n3202 = n2761 & n3201;
  assign n3203 = ~n1186 & n1700;
  assign n3204 = ~n904 & ~n2479;
  assign n3205 = n1479 & ~n3204;
  assign n3206 = n462 & n1900;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n3203 & n3207;
  assign n3209 = pi027 & n1398;
  assign n3210 = pi022 & n1684;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = n3208 & n3211;
  assign n3213 = n623 & n3212;
  assign n3214 = ~n1037 & ~n3191;
  assign n3215 = ~n2057 & ~n2909;
  assign n3216 = n2670 & n3215;
  assign n3217 = n1803 & n3216;
  assign n3218 = ~n3214 & n3217;
  assign n3219 = n3213 & n3218;
  assign n3220 = n3202 & n3219;
  assign n3221 = n3195 & n3220;
  assign n3222 = ~pi019 & n1760;
  assign n3223 = ~pi061 & n638;
  assign n3224 = n717 & n3223;
  assign n3225 = ~n458 & ~n648;
  assign n3226 = n690 & ~n3225;
  assign n3227 = ~pi014 & ~n333;
  assign n3228 = n1949 & n3227;
  assign n3229 = ~n3226 & ~n3228;
  assign n3230 = ~n3224 & n3229;
  assign n3231 = ~n501 & n3230;
  assign n3232 = ~n3222 & n3231;
  assign n3233 = n591 & n1241;
  assign n3234 = n1840 & ~n2121;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = ~n1694 & n3235;
  assign n3237 = ~n782 & ~n2855;
  assign n3238 = ~n319 & n2419;
  assign n3239 = ~pi108 & n1618;
  assign n3240 = n347 & n3239;
  assign n3241 = ~n3238 & ~n3240;
  assign n3242 = n3237 & n3241;
  assign n3243 = n3236 & n3242;
  assign n3244 = ~n643 & ~n1646;
  assign n3245 = ~n844 & n3244;
  assign n3246 = n588 & ~n3245;
  assign n3247 = ~pi074 & n2816;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = n3243 & n3248;
  assign n3250 = n3232 & n3249;
  assign n3251 = pi108 & n2242;
  assign n3252 = n2178 & n2209;
  assign n3253 = ~n3251 & n3252;
  assign n3254 = n2749 & n3253;
  assign n3255 = pi013 & ~n1392;
  assign n3256 = ~n649 & ~n3255;
  assign n3257 = ~n2225 & n3256;
  assign n3258 = n336 & n464;
  assign n3259 = n269 & n1241;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = n3257 & n3260;
  assign n3262 = n1973 & n2088;
  assign n3263 = ~n1101 & ~n3262;
  assign n3264 = ~n2710 & n3263;
  assign n3265 = n686 & n2111;
  assign n3266 = ~n2126 & ~n3265;
  assign n3267 = n234 & ~n3266;
  assign n3268 = n2737 & ~n3267;
  assign n3269 = n3264 & n3268;
  assign n3270 = n3261 & n3269;
  assign n3271 = n3254 & n3270;
  assign n3272 = ~pi022 & ~n2248;
  assign n3273 = pi012 & ~n903;
  assign n3274 = n1969 & n3273;
  assign n3275 = ~pi023 & n572;
  assign n3276 = ~n3274 & ~n3275;
  assign n3277 = n224 & n1422;
  assign n3278 = ~n2778 & ~n3277;
  assign n3279 = n3276 & n3278;
  assign n3280 = ~n3272 & n3279;
  assign n3281 = n3271 & n3280;
  assign n3282 = n3250 & n3281;
  assign n3283 = n1515 & n3282;
  assign n3284 = n3221 & n3283;
  assign po16 = ~n3168 | ~n3284;
  assign n3286 = ~pi015 & n2331;
  assign n3287 = ~n2840 & ~n3151;
  assign n3288 = ~n3286 & n3287;
  assign n3289 = ~pi012 & ~n3288;
  assign n3290 = ~n412 & ~n2459;
  assign n3291 = ~n3289 & n3290;
  assign n3292 = n342 & n561;
  assign n3293 = n225 & n3292;
  assign n3294 = ~n1589 & ~n3293;
  assign n3295 = n1247 & n3294;
  assign n3296 = pi007 & n2866;
  assign n3297 = ~n2532 & ~n3296;
  assign n3298 = n574 & ~n3297;
  assign n3299 = ~n390 & ~n3298;
  assign n3300 = n3295 & n3299;
  assign n3301 = n548 & n867;
  assign n3302 = ~n1868 & ~n3301;
  assign n3303 = ~n464 & ~n2339;
  assign n3304 = n317 & ~n3303;
  assign n3305 = ~n1877 & ~n3304;
  assign n3306 = n3302 & n3305;
  assign n3307 = n3300 & n3306;
  assign n3308 = n3291 & n3307;
  assign n3309 = n499 & ~n911;
  assign n3310 = n1578 & n3309;
  assign n3311 = ~pi013 & n928;
  assign n3312 = n974 & n2159;
  assign n3313 = ~pi014 & ~n2111;
  assign n3314 = ~n2334 & ~n3313;
  assign n3315 = n690 & ~n3314;
  assign n3316 = ~n3312 & ~n3315;
  assign n3317 = ~n3311 & n3316;
  assign n3318 = n3310 & n3317;
  assign n3319 = pi023 & n451;
  assign n3320 = n2926 & ~n3319;
  assign n3321 = n741 & ~n3320;
  assign n3322 = ~pi019 & n3321;
  assign n3323 = n1473 & n2729;
  assign n3324 = ~n1481 & ~n3323;
  assign n3325 = n458 & ~n3324;
  assign n3326 = n392 & n1598;
  assign n3327 = ~n773 & n843;
  assign n3328 = n588 & ~n736;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = n3326 & ~n3329;
  assign n3331 = ~n3325 & ~n3330;
  assign n3332 = ~n3322 & n3331;
  assign n3333 = ~n2576 & ~n2957;
  assign n3334 = n1940 & n3333;
  assign n3335 = ~n1970 & n3334;
  assign n3336 = n3332 & n3335;
  assign n3337 = n3318 & n3336;
  assign n3338 = ~pi074 & n2880;
  assign n3339 = ~n1609 & ~n1993;
  assign n3340 = n784 & n789;
  assign n3341 = ~n791 & ~n3340;
  assign n3342 = ~n512 & n3341;
  assign n3343 = n2333 & ~n3342;
  assign n3344 = pi019 & n467;
  assign n3345 = ~n1153 & ~n1304;
  assign n3346 = ~n3344 & n3345;
  assign n3347 = n2902 & ~n3346;
  assign n3348 = ~n3343 & ~n3347;
  assign n3349 = n3339 & n3348;
  assign n3350 = ~n3338 & n3349;
  assign n3351 = ~n1579 & ~n2501;
  assign n3352 = n432 & ~n3351;
  assign n3353 = n270 & n2585;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = ~n1978 & ~n2746;
  assign n3356 = n815 & ~n3355;
  assign n3357 = ~n2369 & ~n3356;
  assign n3358 = n865 & ~n3357;
  assign n3359 = n1477 & n1950;
  assign n3360 = n1741 & n3009;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3358 & n3361;
  assign n3363 = ~n421 & n3362;
  assign n3364 = n3354 & n3363;
  assign n3365 = n3350 & n3364;
  assign n3366 = n3337 & n3365;
  assign n3367 = n3308 & n3366;
  assign n3368 = ~n1760 & ~n2542;
  assign n3369 = n2188 & n3368;
  assign n3370 = n1085 & n2093;
  assign n3371 = ~n504 & ~n3370;
  assign n3372 = ~n898 & n3371;
  assign n3373 = ~n2487 & n3372;
  assign n3374 = n345 & n2372;
  assign n3375 = ~pi005 & ~n3026;
  assign n3376 = ~n337 & ~n3375;
  assign n3377 = n1847 & ~n3376;
  assign n3378 = ~n2492 & ~n3377;
  assign n3379 = ~n3374 & n3378;
  assign n3380 = ~n1819 & ~n2462;
  assign n3381 = ~n1236 & n3380;
  assign n3382 = n3379 & n3381;
  assign n3383 = n3373 & n3382;
  assign n3384 = pi019 & n2636;
  assign n3385 = ~n357 & n2525;
  assign n3386 = ~pi015 & n2948;
  assign n3387 = pi010 & n3386;
  assign n3388 = ~n3385 & ~n3387;
  assign n3389 = ~n3384 & n3388;
  assign n3390 = n3383 & n3389;
  assign n3391 = n3369 & n3390;
  assign n3392 = n3257 & n3391;
  assign n3393 = n3367 & n3392;
  assign n3394 = n1547 & n2838;
  assign n3395 = ~n2307 & ~n3394;
  assign n3396 = n1833 & n2074;
  assign n3397 = n458 & n2126;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = n3395 & n3398;
  assign n3400 = ~n1401 & n3399;
  assign n3401 = ~n639 & ~n1345;
  assign n3402 = ~n2027 & n3401;
  assign n3403 = n2249 & n3402;
  assign n3404 = n3400 & n3403;
  assign n3405 = ~n1453 & n3404;
  assign n3406 = n636 & n3264;
  assign n3407 = n1833 & n1834;
  assign n3408 = n1090 & n1953;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = ~n1088 & n3409;
  assign n3411 = n342 & n2259;
  assign n3412 = n483 & n1664;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~pi014 & n702;
  assign n3415 = n892 & n3414;
  assign n3416 = ~n1893 & ~n2629;
  assign n3417 = n517 & ~n3416;
  assign n3418 = ~n3415 & ~n3417;
  assign n3419 = n3413 & n3418;
  assign n3420 = n3410 & n3419;
  assign n3421 = n1557 & n3420;
  assign n3422 = ~n955 & n3421;
  assign n3423 = n3406 & n3422;
  assign n3424 = n2979 & n3423;
  assign n3425 = n1311 & n3424;
  assign n3426 = n3405 & n3425;
  assign n3427 = n3393 & n3426;
  assign n3428 = ~n667 & n3164;
  assign n3429 = n609 & n1154;
  assign n3430 = ~n1141 & ~n1582;
  assign n3431 = ~n3429 & n3430;
  assign n3432 = n613 & ~n1140;
  assign n3433 = ~pi022 & n1825;
  assign n3434 = n1126 & n1878;
  assign n3435 = ~n3433 & ~n3434;
  assign n3436 = n541 & ~n3435;
  assign n3437 = n471 & n1619;
  assign n3438 = n836 & n3437;
  assign n3439 = ~n3436 & ~n3438;
  assign n3440 = n3432 & n3439;
  assign n3441 = n3431 & n3440;
  assign n3442 = ~n383 & ~n3441;
  assign n3443 = n876 & n3033;
  assign n3444 = ~n2228 & ~n2271;
  assign n3445 = pi018 & ~n3444;
  assign n3446 = ~n1277 & ~n3445;
  assign n3447 = ~n374 & n375;
  assign n3448 = ~n3446 & n3447;
  assign n3449 = n1733 & ~n3448;
  assign n3450 = n3443 & n3449;
  assign n3451 = ~n3442 & n3450;
  assign n3452 = n2420 & ~n3277;
  assign n3453 = ~n1892 & n3452;
  assign n3454 = ~pi018 & n2512;
  assign n3455 = ~n732 & ~n1607;
  assign n3456 = n678 & ~n3455;
  assign n3457 = ~n3454 & ~n3456;
  assign n3458 = n710 & n2845;
  assign n3459 = pi012 & n712;
  assign n3460 = ~n3458 & ~n3459;
  assign n3461 = ~pi015 & ~n3460;
  assign n3462 = ~n559 & ~n572;
  assign n3463 = pi023 & ~n3462;
  assign n3464 = ~n3461 & ~n3463;
  assign n3465 = n3457 & n3464;
  assign n3466 = n1805 & n3465;
  assign n3467 = n3453 & n3466;
  assign n3468 = n3451 & n3467;
  assign n3469 = n3428 & n3468;
  assign n3470 = n3427 & n3469;
  assign n3471 = n3221 & n3470;
  assign po17 = ~n1524 | ~n3471;
  assign n3473 = ~n634 & ~n2931;
  assign n3474 = ~n427 & ~n3370;
  assign n3475 = ~n229 & ~n342;
  assign n3476 = n1848 & ~n3475;
  assign n3477 = n3474 & ~n3476;
  assign n3478 = n3473 & n3477;
  assign n3479 = pi003 & n1246;
  assign n3480 = ~n3224 & ~n3479;
  assign n3481 = n482 & n1303;
  assign n3482 = ~pi021 & n751;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = n3480 & n3483;
  assign n3485 = n3478 & n3484;
  assign po18 = ~n3452 | ~n3485;
  assign n3487 = n1273 & n2590;
  assign n3488 = n3077 & n3487;
  assign n3489 = ~n2563 & n2899;
  assign n3490 = n1616 & n3024;
  assign n3491 = n3489 & n3490;
  assign n3492 = n3488 & n3491;
  assign n3493 = n511 & n937;
  assign n3494 = ~pi013 & n3493;
  assign n3495 = n2425 & ~n3494;
  assign n3496 = n233 & n2159;
  assign n3497 = pi013 & n2251;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = n2925 & n3498;
  assign n3500 = n480 & n494;
  assign n3501 = n399 & n561;
  assign n3502 = ~n2180 & ~n3501;
  assign n3503 = ~n3292 & n3502;
  assign n3504 = ~n3500 & n3503;
  assign n3505 = pi002 & ~n3504;
  assign n3506 = ~n397 & n3460;
  assign n3507 = ~n3505 & n3506;
  assign n3508 = n3499 & n3507;
  assign n3509 = ~n1236 & ~n1298;
  assign n3510 = n2361 & n3509;
  assign n3511 = n984 & n1291;
  assign n3512 = ~n2269 & ~n3511;
  assign n3513 = ~n2408 & n3512;
  assign n3514 = n3510 & n3513;
  assign n3515 = n3508 & n3514;
  assign n3516 = n3495 & n3515;
  assign n3517 = ~n2257 & n3516;
  assign n3518 = n3492 & n3517;
  assign n3519 = n1081 & n1642;
  assign n3520 = ~n1453 & n3519;
  assign n3521 = ~n511 & ~n1735;
  assign n3522 = ~n786 & n3521;
  assign n3523 = n701 & ~n3522;
  assign n3524 = n451 & n735;
  assign n3525 = ~n267 & n3524;
  assign n3526 = ~n869 & ~n3525;
  assign n3527 = n2524 & n3526;
  assign n3528 = n2968 & n3527;
  assign n3529 = ~n3523 & n3528;
  assign n3530 = n3520 & n3529;
  assign n3531 = n3140 & n3530;
  assign n3532 = n3518 & n3531;
  assign n3533 = n2464 & n2631;
  assign n3534 = ~n2062 & n3533;
  assign n3535 = ~n867 & n3534;
  assign n3536 = n2964 & n3535;
  assign n3537 = ~n2346 & n3536;
  assign n3538 = ~n911 & n3537;
  assign n3539 = ~n3151 & n3538;
  assign n3540 = n2460 & n2837;
  assign n3541 = ~n1222 & ~n1398;
  assign n3542 = ~n1793 & n3401;
  assign n3543 = n3084 & n3542;
  assign n3544 = n3541 & n3543;
  assign n3545 = ~pi027 & ~n2025;
  assign n3546 = ~n2696 & ~n3545;
  assign n3547 = n2217 & n3546;
  assign n3548 = n3544 & n3547;
  assign n3549 = ~n630 & ~n1112;
  assign n3550 = ~n1070 & ~n3549;
  assign n3551 = pi022 & n1293;
  assign n3552 = n483 & n659;
  assign n3553 = ~n3551 & ~n3552;
  assign n3554 = ~pi013 & n1291;
  assign n3555 = pi014 & n3554;
  assign n3556 = n3553 & ~n3555;
  assign n3557 = ~n634 & n3556;
  assign n3558 = ~n383 & n1004;
  assign n3559 = n443 & n1827;
  assign n3560 = ~n2097 & ~n3559;
  assign n3561 = ~n486 & ~n2768;
  assign n3562 = n3560 & n3561;
  assign n3563 = n2037 & n3562;
  assign n3564 = ~n3558 & n3563;
  assign n3565 = n3557 & n3564;
  assign n3566 = ~n3550 & n3565;
  assign n3567 = n3548 & n3566;
  assign n3568 = n2157 & n3049;
  assign n3569 = n3567 & n3568;
  assign n3570 = n3540 & n3569;
  assign n3571 = n3539 & n3570;
  assign po19 = ~n3532 | ~n3571;
  assign n3573 = n1274 & n2294;
  assign n3574 = pi011 & n2111;
  assign n3575 = n3135 & n3574;
  assign n3576 = ~n1047 & ~n3511;
  assign n3577 = n2420 & ~n2549;
  assign n3578 = n3127 & n3577;
  assign n3579 = n3576 & n3578;
  assign n3580 = ~n3575 & n3579;
  assign n3581 = n3573 & n3580;
  assign n3582 = ~n705 & n906;
  assign n3583 = ~n2329 & ~n2498;
  assign n3584 = ~n3582 & n3583;
  assign n3585 = n802 & ~n3131;
  assign n3586 = n815 & n2444;
  assign n3587 = ~n3585 & ~n3586;
  assign n3588 = ~n3019 & ~n3118;
  assign n3589 = n3587 & n3588;
  assign n3590 = n3584 & n3589;
  assign n3591 = ~n2589 & n3590;
  assign n3592 = pi014 & n2252;
  assign n3593 = n3591 & ~n3592;
  assign n3594 = n2807 & n3593;
  assign n3595 = n3581 & n3594;
  assign po20 = ~n3570 | ~n3595;
  assign n3597 = n1699 & ~n3558;
  assign n3598 = n3020 & n3597;
  assign n3599 = ~n2943 & n3147;
  assign n3600 = pi027 & n2023;
  assign n3601 = n1072 & n2200;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = n3599 & n3602;
  assign n3604 = n3598 & n3603;
  assign n3605 = n777 & n1703;
  assign n3606 = ~pi009 & n3605;
  assign n3607 = ~n1260 & ~n3606;
  assign n3608 = ~n2174 & n3607;
  assign n3609 = ~n2205 & n3608;
  assign n3610 = ~n916 & n3609;
  assign n3611 = ~n1801 & n3584;
  assign n3612 = n3610 & n3611;
  assign n3613 = ~n789 & n903;
  assign n3614 = ~n1876 & ~n2288;
  assign n3615 = ~n3613 & n3614;
  assign n3616 = n1262 & ~n3615;
  assign n3617 = ~n2317 & ~n3616;
  assign n3618 = ~n1901 & n3617;
  assign n3619 = n3612 & n3618;
  assign n3620 = n346 & n659;
  assign n3621 = n450 & n663;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = ~n383 & ~n3622;
  assign n3624 = ~n1871 & ~n3623;
  assign n3625 = n3038 & n3624;
  assign n3626 = ~n2163 & n3625;
  assign n3627 = n3619 & n3626;
  assign n3628 = n3604 & n3627;
  assign n3629 = n318 & ~n3190;
  assign n3630 = ~n345 & n1243;
  assign n3631 = n1848 & ~n3630;
  assign n3632 = ~n3629 & ~n3631;
  assign n3633 = ~n1885 & n3632;
  assign n3634 = n382 & n1884;
  assign n3635 = ~n1314 & ~n3634;
  assign n3636 = n3633 & n3635;
  assign n3637 = n1587 & n3636;
  assign n3638 = ~n493 & n3637;
  assign n3639 = n2295 & n3638;
  assign n3640 = pi011 & n2177;
  assign n3641 = n234 & n1259;
  assign n3642 = ~n1902 & ~n3641;
  assign n3643 = ~n3640 & n3642;
  assign n3644 = ~n234 & n1904;
  assign n3645 = ~n894 & ~n2186;
  assign n3646 = ~n3644 & n3645;
  assign n3647 = n3643 & n3646;
  assign n3648 = ~n1701 & n3647;
  assign n3649 = ~n2403 & ~n3135;
  assign n3650 = n3574 & ~n3649;
  assign n3651 = ~n2252 & ~n3585;
  assign n3652 = ~n890 & n3651;
  assign n3653 = ~n3650 & n3652;
  assign n3654 = n3648 & n3653;
  assign n3655 = ~n2007 & ~n2207;
  assign n3656 = n3654 & n3655;
  assign n3657 = n3639 & n3656;
  assign n3658 = n3628 & n3657;
  assign n3659 = ~n302 & n1029;
  assign n3660 = ~n1015 & ~n3659;
  assign n3661 = ~n356 & n1024;
  assign n3662 = n3660 & n3661;
  assign n3663 = n3171 & ~n3177;
  assign n3664 = n3662 & ~n3663;
  assign n3665 = ~n3193 & n3664;
  assign n3666 = n3188 & n3665;
  assign n3667 = n1997 & n3666;
  assign n3668 = n3658 & n3667;
  assign n3669 = n953 & n3528;
  assign n3670 = n457 & n1763;
  assign n3671 = n3489 & n3670;
  assign n3672 = n3669 & n3671;
  assign n3673 = ~n551 & ~n588;
  assign n3674 = n3433 & ~n3673;
  assign n3675 = ~n2752 & ~n3674;
  assign n3676 = ~n1130 & n1862;
  assign n3677 = n3675 & ~n3676;
  assign n3678 = n502 & n632;
  assign n3679 = ~n1726 & ~n3678;
  assign n3680 = ~n383 & ~n3679;
  assign n3681 = ~n273 & n551;
  assign n3682 = n1643 & n3681;
  assign n3683 = n985 & n1833;
  assign n3684 = ~n2112 & ~n3683;
  assign n3685 = ~n1282 & n3684;
  assign n3686 = ~n3682 & n3685;
  assign n3687 = ~n3680 & n3686;
  assign n3688 = n3473 & n3687;
  assign n3689 = n3677 & n3688;
  assign n3690 = n2811 & n3261;
  assign n3691 = n3689 & n3690;
  assign n3692 = n2588 & n3691;
  assign n3693 = n3672 & n3692;
  assign n3694 = ~n2020 & ~n2024;
  assign n3695 = pi027 & ~n3694;
  assign n3696 = ~n3162 & ~n3695;
  assign n3697 = n1748 & n3414;
  assign n3698 = ~n2797 & ~n3697;
  assign n3699 = ~n766 & ~n3698;
  assign n3700 = ~n2688 & ~n3699;
  assign n3701 = ~pi060 & n3021;
  assign n3702 = n1734 & n1735;
  assign n3703 = pi069 & n3702;
  assign n3704 = ~n824 & ~n3703;
  assign n3705 = ~n3701 & n3704;
  assign n3706 = n3700 & n3705;
  assign n3707 = n3696 & n3706;
  assign n3708 = n1105 & n3707;
  assign n3709 = n3202 & n3708;
  assign n3710 = ~n1544 & n1820;
  assign n3711 = ~n1541 & n3710;
  assign n3712 = n1148 & n3711;
  assign n3713 = n3404 & n3712;
  assign n3714 = n311 & n1031;
  assign n3715 = n1033 & n3714;
  assign n3716 = ~n3191 & ~n3715;
  assign n3717 = n3453 & ~n3716;
  assign n3718 = n3713 & n3717;
  assign n3719 = n3709 & n3718;
  assign n3720 = n3693 & n3719;
  assign n3721 = n3668 & n3720;
  assign n3722 = n1530 & n1688;
  assign n3723 = n3106 & n3722;
  assign po21 = ~n3721 | ~n3723;
  assign n3725 = ~n1036 & ~n3191;
  assign n3726 = ~n3199 & ~n3725;
  assign n3727 = ~n287 & n3726;
  assign po22 = ~n3666 | ~n3727;
  assign n3729 = n2017 & n3609;
  assign n3730 = n790 & n2469;
  assign n3731 = ~n2847 & ~n3730;
  assign n3732 = n910 & n934;
  assign n3733 = ~n3100 & ~n3732;
  assign n3734 = ~n2347 & n3733;
  assign n3735 = n3731 & n3734;
  assign n3736 = n1898 & ~n3458;
  assign n3737 = ~n1816 & n3736;
  assign n3738 = ~n810 & n3737;
  assign n3739 = n1330 & n3738;
  assign n3740 = n3735 & n3739;
  assign n3741 = ~n1272 & n3512;
  assign n3742 = pi015 & n3459;
  assign n3743 = ~n703 & ~n3742;
  assign n3744 = n3700 & n3743;
  assign n3745 = n3741 & n3744;
  assign n3746 = n3740 & n3745;
  assign n3747 = n3729 & n3746;
  assign n3748 = ~n333 & n911;
  assign n3749 = ~n1700 & ~n3748;
  assign n3750 = ~n334 & ~n3749;
  assign n3751 = ~n3041 & ~n3750;
  assign n3752 = ~n1264 & ~n2446;
  assign n3753 = n3647 & n3752;
  assign n3754 = ~pi027 & n3555;
  assign n3755 = n3536 & ~n3754;
  assign n3756 = n3753 & n3755;
  assign n3757 = n3751 & n3756;
  assign n3758 = n3747 & n3757;
  assign po23 = ~n3158 | ~n3758;
  assign n3760 = ~pi020 & ~pi122;
  assign n3761 = n223 & ~n3760;
  assign n3762 = n395 & ~n3761;
  assign n3763 = ~n2257 & ~n3762;
  assign n3764 = n1847 & ~n3630;
  assign n3765 = n3763 & ~n3764;
  assign n3766 = n2026 & n3765;
  assign n3767 = n1121 & n3766;
  assign n3768 = ~n1321 & ~n1787;
  assign n3769 = ~n1147 & n3768;
  assign n3770 = ~n622 & n1214;
  assign n3771 = ~n1270 & n3770;
  assign n3772 = n3541 & n3771;
  assign n3773 = n3769 & n3772;
  assign n3774 = n2760 & n3773;
  assign n3775 = n3767 & n3774;
  assign n3776 = pi056 & ~pi122;
  assign n3777 = ~n1164 & ~n3776;
  assign n3778 = n1343 & n3777;
  assign n3779 = n2424 & ~n2894;
  assign n3780 = n1175 & ~n2207;
  assign n3781 = n3779 & n3780;
  assign n3782 = ~n3778 & n3781;
  assign n3783 = ~pi027 & ~n3553;
  assign n3784 = n354 & n1046;
  assign n3785 = n3069 & ~n3784;
  assign n3786 = ~n2419 & n3785;
  assign n3787 = ~n3783 & n3786;
  assign n3788 = n3040 & n3787;
  assign n3789 = n3782 & n3788;
  assign n3790 = n1963 & n2456;
  assign n3791 = n3789 & n3790;
  assign n3792 = n3775 & n3791;
  assign n3793 = ~n1047 & n1238;
  assign n3794 = n1311 & n3793;
  assign n3795 = n2836 & n3405;
  assign n3796 = n3794 & n3795;
  assign n3797 = n1520 & n3099;
  assign n3798 = n3796 & n3797;
  assign n3799 = n3792 & n3798;
  assign n3800 = n1690 & n3693;
  assign po24 = ~n3799 | ~n3800;
  assign n3802 = pi027 & ~n3556;
  assign n3803 = n377 & n1331;
  assign n3804 = ~n3021 & ~n3803;
  assign n3805 = n3624 & n3804;
  assign n3806 = ~n3802 & n3805;
  assign n3807 = ~pi014 & n3554;
  assign n3808 = ~n3162 & ~n3807;
  assign n3809 = ~n614 & n3808;
  assign n3810 = n2679 & n3809;
  assign po25 = ~n3806 | ~n3810;
  assign po26 = n421 | ~n2287;
  assign n3813 = n530 & n1317;
  assign n3814 = n284 & n1421;
  assign n3815 = n258 & n3814;
  assign n3816 = ~n3813 & ~n3815;
  assign n3817 = ~pi056 & n1313;
  assign n3818 = ~n1168 & n1177;
  assign n3819 = n530 & ~n3818;
  assign n3820 = ~n3817 & ~n3819;
  assign n3821 = n3816 & n3820;
  assign n3822 = ~n1347 & ~n1466;
  assign n3823 = n2123 & n3822;
  assign n3824 = ~n1211 & n3823;
  assign n3825 = n1010 & n3824;
  assign n3826 = ~pi045 & ~n3825;
  assign n3827 = ~pi045 & n343;
  assign n3828 = ~pi007 & n290;
  assign n3829 = ~n1470 & ~n3828;
  assign n3830 = n1431 & n3829;
  assign n3831 = n284 & ~n3830;
  assign n3832 = n1669 & ~n3831;
  assign n3833 = n3827 & ~n3832;
  assign n3834 = ~n1320 & ~n1475;
  assign n3835 = n1337 & n3834;
  assign n3836 = n1059 & ~n3835;
  assign n3837 = pi023 & ~n3351;
  assign n3838 = ~n1670 & ~n3837;
  assign n3839 = n3827 & ~n3838;
  assign n3840 = ~pi045 & n439;
  assign n3841 = n337 & n3840;
  assign n3842 = ~n3839 & ~n3841;
  assign n3843 = n1059 & ~n1433;
  assign n3844 = n1062 & ~n3843;
  assign n3845 = ~pi045 & n405;
  assign n3846 = ~n477 & ~n1249;
  assign n3847 = n3845 & ~n3846;
  assign n3848 = ~pi045 & n269;
  assign n3849 = n228 & n3848;
  assign n3850 = ~n3847 & ~n3849;
  assign n3851 = n3844 & n3850;
  assign n3852 = n3842 & n3851;
  assign n3853 = n651 & n1059;
  assign n3854 = ~pi045 & ~n1189;
  assign n3855 = n581 & n3854;
  assign n3856 = ~pi045 & n345;
  assign n3857 = n1341 & n3856;
  assign n3858 = ~n532 & ~n3857;
  assign n3859 = ~n3855 & n3858;
  assign n3860 = ~n3853 & n3859;
  assign n3861 = n3852 & n3860;
  assign n3862 = ~n3836 & n3861;
  assign n3863 = ~n3833 & n3862;
  assign n3864 = ~n3826 & n3863;
  assign n3865 = n3821 & n3864;
  assign n3866 = n2239 & n3865;
  assign n3867 = n1103 & n1616;
  assign n3868 = ~n1286 & n1449;
  assign n3869 = ~n1075 & n1650;
  assign n3870 = n3868 & n3869;
  assign n3871 = n342 & n1631;
  assign n3872 = ~n1679 & ~n3871;
  assign n3873 = ~n1245 & n3872;
  assign n3874 = n1144 & n3873;
  assign n3875 = ~n3429 & n3874;
  assign n3876 = ~n1673 & n3875;
  assign n3877 = ~n382 & ~n1930;
  assign n3878 = ~n3876 & n3877;
  assign n3879 = ~n2045 & ~n3878;
  assign n3880 = n1240 & n3879;
  assign n3881 = n3870 & n3880;
  assign n3882 = n407 & n2056;
  assign n3883 = ~pi003 & ~pi005;
  assign n3884 = n1082 & n3883;
  assign n3885 = ~n3882 & ~n3884;
  assign n3886 = pi005 & pi007;
  assign n3887 = n3871 & ~n3886;
  assign n3888 = n574 & n3025;
  assign n3889 = n345 & n1769;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = ~n3887 & n3890;
  assign n3892 = n3885 & n3891;
  assign n3893 = ~n1673 & n3892;
  assign n3894 = n1930 & ~n3893;
  assign n3895 = ~n1747 & ~n3894;
  assign n3896 = n3881 & n3895;
  assign n3897 = n3867 & n3896;
  assign n3898 = n1123 & ~n1129;
  assign n3899 = n3432 & ~n3898;
  assign n3900 = ~n544 & ~n1651;
  assign n3901 = ~n1125 & n3900;
  assign n3902 = n3899 & n3901;
  assign n3903 = n284 & n1063;
  assign n3904 = n574 & n3903;
  assign n3905 = n1114 & ~n1705;
  assign n3906 = ~n1066 & n3905;
  assign n3907 = n284 & ~n3906;
  assign n3908 = ~n1134 & ~n1676;
  assign n3909 = ~n3907 & n3908;
  assign n3910 = ~n3904 & n3909;
  assign n3911 = n392 & ~n1216;
  assign n3912 = ~n1283 & ~n3911;
  assign n3913 = n609 & ~n3912;
  assign n3914 = n399 & n1631;
  assign n3915 = ~n1118 & ~n3914;
  assign n3916 = ~n3913 & n3915;
  assign n3917 = ~n1087 & ~n1678;
  assign n3918 = n3916 & n3917;
  assign n3919 = n3910 & n3918;
  assign n3920 = n3902 & n3919;
  assign n3921 = ~n383 & ~n3920;
  assign n3922 = ~n1280 & n2058;
  assign n3923 = ~n2220 & n3922;
  assign n3924 = ~n3921 & n3923;
  assign n3925 = n3897 & n3924;
  assign n3926 = ~pi039 & ~n3925;
  assign n3927 = n1728 & ~n1744;
  assign n3928 = ~n1915 & n1936;
  assign n3929 = n3927 & ~n3928;
  assign n3930 = pi108 & ~n1739;
  assign n3931 = ~pi122 & n3930;
  assign n3932 = ~pi039 & n1928;
  assign n3933 = ~n1918 & ~n3932;
  assign n3934 = ~n1930 & ~n3933;
  assign n3935 = ~n3931 & n3934;
  assign n3936 = ~n3929 & ~n3935;
  assign n3937 = ~pi056 & ~pi122;
  assign n3938 = n258 & ~n3173;
  assign n3939 = ~pi045 & n258;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = ~n3937 & n3940;
  assign n3942 = ~n1038 & ~n3941;
  assign n3943 = ~pi056 & n230;
  assign n3944 = ~pi045 & n337;
  assign n3945 = ~n3943 & ~n3944;
  assign n3946 = n297 & ~n3945;
  assign n3947 = ~n3182 & n3937;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = ~n3172 & ~n3940;
  assign n3950 = n3948 & ~n3949;
  assign n3951 = ~pi056 & ~n3184;
  assign n3952 = n3950 & ~n3951;
  assign n3953 = ~n3942 & n3952;
  assign n3954 = ~n2668 & n3953;
  assign n3955 = n3936 & n3954;
  assign n3956 = ~n3926 & n3955;
  assign n3957 = pi011 & n3121;
  assign n3958 = n777 & n1734;
  assign n3959 = ~n1787 & ~n3958;
  assign n3960 = ~n3957 & n3959;
  assign n3961 = n3956 & n3960;
  assign n3962 = n3866 & n3961;
  assign n3963 = n1696 & ~n2537;
  assign n3964 = ~n2778 & n3963;
  assign n3965 = n3793 & n3964;
  assign n3966 = n224 & n1565;
  assign n3967 = ~n390 & ~n3966;
  assign n3968 = n1587 & n3967;
  assign n3969 = ~n1574 & ~n1588;
  assign n3970 = ~n1534 & n3969;
  assign n3971 = n269 & n496;
  assign n3972 = n3970 & ~n3971;
  assign n3973 = ~n383 & ~n3972;
  assign n3974 = ~n1965 & ~n3973;
  assign n3975 = n3710 & n3974;
  assign n3976 = n3968 & n3975;
  assign n3977 = n3965 & n3976;
  assign n3978 = ~pi039 & ~n3977;
  assign n3979 = n234 & n1902;
  assign n3980 = ~pi011 & n3979;
  assign n3981 = ~n2275 & ~n3980;
  assign n3982 = ~n1528 & n3845;
  assign n3983 = ~pi045 & n982;
  assign n3984 = pi015 & pi122;
  assign n3985 = n3983 & ~n3984;
  assign n3986 = n789 & n3985;
  assign n3987 = ~n3982 & ~n3986;
  assign n3988 = n3981 & n3987;
  assign n3989 = pi034 & ~pi039;
  assign n3990 = n2095 & n3989;
  assign n3991 = ~n2215 & ~n3990;
  assign n3992 = n1267 & n3845;
  assign n3993 = ~pi022 & n3992;
  assign n3994 = ~pi011 & n2910;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = n3991 & n3995;
  assign n3997 = n3988 & n3996;
  assign n3998 = n802 & n2298;
  assign n3999 = n232 & n1930;
  assign n4000 = ~n1835 & ~n1875;
  assign n4001 = n3999 & ~n4000;
  assign n4002 = ~n3198 & ~n4001;
  assign n4003 = ~n3998 & n4002;
  assign n4004 = pi023 & pi039;
  assign n4005 = n569 & ~n4004;
  assign n4006 = ~n855 & ~n4005;
  assign n4007 = n1217 & ~n4006;
  assign n4008 = ~n475 & n3845;
  assign n4009 = ~pi039 & n575;
  assign n4010 = ~pi045 & n4009;
  assign n4011 = ~n4008 & ~n4010;
  assign n4012 = ~n4007 & n4011;
  assign n4013 = n3200 & n4012;
  assign n4014 = n4003 & n4013;
  assign n4015 = n1274 & n4014;
  assign n4016 = n3997 & n4015;
  assign n4017 = ~n1423 & n1930;
  assign n4018 = n2667 & ~n4017;
  assign n4019 = n4016 & n4018;
  assign n4020 = ~n3978 & n4019;
  assign n4021 = ~n1706 & n1758;
  assign n4022 = n1185 & n1969;
  assign n4023 = n284 & n633;
  assign n4024 = n764 & n872;
  assign n4025 = ~pi039 & n551;
  assign n4026 = n2801 & n4025;
  assign n4027 = ~n4024 & ~n4026;
  assign n4028 = ~n4023 & n4027;
  assign n4029 = ~n4022 & n4028;
  assign n4030 = n4021 & n4029;
  assign n4031 = ~pi001 & n941;
  assign n4032 = n3608 & ~n4031;
  assign n4033 = n2314 & n4032;
  assign n4034 = n4030 & n4033;
  assign n4035 = ~pi004 & ~pi108;
  assign n4036 = n2316 & ~n4035;
  assign n4037 = n444 & n1619;
  assign n4038 = ~n830 & ~n4037;
  assign n4039 = ~n4036 & n4038;
  assign n4040 = ~pi010 & n1749;
  assign n4041 = ~n893 & ~n1900;
  assign n4042 = n903 & ~n4041;
  assign n4043 = n354 & n1199;
  assign n4044 = n268 & n4043;
  assign n4045 = ~n4042 & ~n4044;
  assign n4046 = ~n4040 & n4045;
  assign n4047 = ~n1700 & n4046;
  assign n4048 = n4039 & n4047;
  assign n4049 = n4034 & n4048;
  assign n4050 = ~n1974 & ~n2204;
  assign n4051 = n334 & ~n4050;
  assign n4052 = n1208 & n3110;
  assign n4053 = ~n3620 & ~n4052;
  assign n4054 = ~pi045 & ~n4053;
  assign n4055 = pi011 & ~n547;
  assign n4056 = ~n2296 & n4055;
  assign n4057 = ~n4054 & ~n4056;
  assign n4058 = ~n4051 & n4057;
  assign n4059 = n4049 & n4058;
  assign n4060 = n4020 & n4059;
  assign n4061 = n3168 & n4060;
  assign po28 = ~n3962 | ~n4061;
  assign n4063 = n942 & n3495;
  assign n4064 = n734 & ~n749;
  assign n4065 = ~n2270 & ~n4064;
  assign n4066 = n482 & ~n4065;
  assign n4067 = n735 & n1536;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n387 & ~n2586;
  assign n4070 = n376 & n468;
  assign n4071 = ~n1826 & ~n4070;
  assign n4072 = n384 & ~n4071;
  assign n4073 = n230 & n1278;
  assign n4074 = pi020 & n394;
  assign n4075 = ~n2304 & n4074;
  assign n4076 = ~n4073 & ~n4075;
  assign n4077 = n1126 & ~n4076;
  assign n4078 = ~n4072 & ~n4077;
  assign n4079 = ~n4069 & n4078;
  assign n4080 = n4068 & n4079;
  assign n4081 = ~n1879 & ~n3990;
  assign n4082 = n4080 & n4081;
  assign n4083 = n4063 & n4082;
  assign n4084 = ~n683 & ~n2264;
  assign n4085 = n3520 & ~n4084;
  assign n4086 = n1593 & n4085;
  assign n4087 = n3794 & n4086;
  assign n4088 = ~n1661 & n4087;
  assign n4089 = ~pi039 & ~n4088;
  assign n4090 = n3672 & ~n4089;
  assign n4091 = n4083 & n4090;
  assign n4092 = ~n939 & n2322;
  assign n4093 = n701 & n926;
  assign n4094 = n458 & n4093;
  assign n4095 = ~n2175 & ~n3090;
  assign n4096 = ~n4094 & n4095;
  assign n4097 = n3766 & n4096;
  assign n4098 = n2218 & n4097;
  assign n4099 = n4092 & n4098;
  assign n4100 = pi001 & ~pi002;
  assign n4101 = pi000 & n1372;
  assign n4102 = n4100 & n4101;
  assign n4103 = n619 & n4102;
  assign n4104 = n225 & n2143;
  assign n4105 = pi000 & ~n4104;
  assign n4106 = n1372 & ~n4105;
  assign n4107 = n225 & n4101;
  assign n4108 = n274 & n4107;
  assign n4109 = n343 & n4108;
  assign n4110 = ~pi017 & n752;
  assign n4111 = n4109 & n4110;
  assign n4112 = pi016 & n4111;
  assign n4113 = ~n4106 & ~n4112;
  assign n4114 = n717 & ~n4113;
  assign n4115 = n251 & n4108;
  assign n4116 = n289 & n4101;
  assign n4117 = n592 & n4116;
  assign n4118 = n317 & n4117;
  assign n4119 = ~n4115 & ~n4118;
  assign n4120 = n1728 & ~n4119;
  assign n4121 = ~n4114 & ~n4120;
  assign n4122 = ~n4103 & n4121;
  assign n4123 = n346 & n4117;
  assign n4124 = n415 & n4116;
  assign n4125 = pi008 & n4124;
  assign n4126 = ~n654 & n1369;
  assign n4127 = ~n2629 & ~n4126;
  assign n4128 = n4125 & ~n4127;
  assign n4129 = ~n4123 & ~n4128;
  assign n4130 = ~pi008 & n4124;
  assign n4131 = pi010 & pi011;
  assign n4132 = pi009 & ~n4131;
  assign n4133 = n4130 & n4132;
  assign n4134 = n4129 & ~n4133;
  assign n4135 = n354 & ~n4134;
  assign n4136 = ~n4108 & ~n4117;
  assign n4137 = ~pi004 & ~n4136;
  assign n4138 = pi016 & ~n1414;
  assign n4139 = ~n1499 & n4138;
  assign n4140 = n4109 & ~n4139;
  assign n4141 = pi002 & ~n1630;
  assign n4142 = n4101 & ~n4141;
  assign n4143 = pi001 & pi006;
  assign n4144 = ~n268 & n4143;
  assign n4145 = ~n2143 & n4107;
  assign n4146 = ~n4144 & n4145;
  assign n4147 = ~n4142 & ~n4146;
  assign n4148 = ~n4140 & n4147;
  assign n4149 = ~n4137 & n4148;
  assign n4150 = n354 & ~n4149;
  assign n4151 = ~pi056 & n4150;
  assign n4152 = ~n4135 & ~n4151;
  assign n4153 = n4122 & n4152;
  assign n4154 = n3071 & n4153;
  assign n4155 = n4099 & n4154;
  assign n4156 = n4091 & n4155;
  assign n4157 = n909 & n2845;
  assign n4158 = pi010 & n4157;
  assign n4159 = n3539 & ~n4158;
  assign n4160 = ~n703 & ~n3958;
  assign n4161 = ~n458 & ~n4160;
  assign n4162 = ~n3732 & ~n3742;
  assign n4163 = n579 & n767;
  assign n4164 = ~pi007 & n234;
  assign n4165 = n974 & ~n4164;
  assign n4166 = ~n791 & ~n1735;
  assign n4167 = pi007 & ~n4166;
  assign n4168 = ~n2288 & ~n4167;
  assign n4169 = ~n4165 & n4168;
  assign n4170 = n4163 & ~n4169;
  assign n4171 = ~n3109 & ~n4170;
  assign n4172 = n4162 & n4171;
  assign n4173 = n3654 & n4172;
  assign n4174 = n3144 & n4173;
  assign n4175 = ~n4161 & n4174;
  assign n4176 = n4159 & n4175;
  assign n4177 = n659 & n3827;
  assign n4178 = pi022 & n3992;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = n934 & n2204;
  assign n4181 = ~n3606 & ~n4180;
  assign n4182 = n2912 & n4181;
  assign n4183 = n3395 & n4182;
  assign n4184 = n4179 & n4183;
  assign n4185 = n1789 & n3200;
  assign n4186 = n413 & n4185;
  assign n4187 = n4184 & n4186;
  assign n4188 = n3130 & n4187;
  assign n4189 = n3428 & n4188;
  assign n4190 = n4176 & n4189;
  assign n4191 = n4156 & n4190;
  assign po29 = ~n3956 | ~n4191;
  assign n4193 = n1423 & ~n4052;
  assign n4194 = ~pi045 & ~n4193;
  assign n4195 = ~n2678 & ~n4194;
  assign n4196 = ~n1914 & ~n4195;
  assign n4197 = n3414 & n3877;
  assign n4198 = ~pi045 & n1478;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = n1208 & ~n4199;
  assign n4201 = ~n458 & ~n863;
  assign n4202 = n1914 & ~n4201;
  assign n4203 = n983 & n4202;
  assign n4204 = ~n1529 & n4012;
  assign n4205 = ~n4203 & n4204;
  assign n4206 = ~n4200 & n4205;
  assign n4207 = ~n4196 & n4206;
  assign n4208 = n4002 & n4207;
  assign n4209 = n3865 & n4208;
  assign n4210 = ~n382 & n472;
  assign n4211 = ~pi045 & n375;
  assign n4212 = pi019 & n1930;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = ~n4210 & n4213;
  assign n4215 = n450 & ~n4214;
  assign n4216 = n662 & n4215;
  assign n4217 = n659 & n3856;
  assign n4218 = pi122 & n4217;
  assign n4219 = n3620 & n3877;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = ~n4177 & n4220;
  assign n4222 = ~n4216 & n4221;
  assign n4223 = ~n1848 & n4222;
  assign n4224 = n2420 & n4223;
  assign n4225 = ~n1301 & ~n1306;
  assign n4226 = n480 & n1299;
  assign n4227 = ~pi007 & n4226;
  assign n4228 = n4225 & ~n4227;
  assign n4229 = n2503 & n4228;
  assign n4230 = n383 & ~n446;
  assign n4231 = n1639 & ~n4230;
  assign n4232 = n2264 & ~n4231;
  assign n4233 = n4229 & n4232;
  assign n4234 = ~n3481 & n4233;
  assign n4235 = ~pi039 & ~n4234;
  assign n4236 = pi019 & ~n457;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = n4224 & n4237;
  assign n4239 = n4153 & n4238;
  assign po30 = ~n4209 | ~n4239;
  assign n4241 = n557 & n2513;
  assign n4242 = n1876 & n4163;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = ~n4157 & n4243;
  assign n4245 = ~n381 & n4244;
  assign n4246 = ~n984 & n2468;
  assign n4247 = ~n917 & ~n4246;
  assign n4248 = n2896 & n4247;
  assign n4249 = n4245 & n4248;
  assign n4250 = n2425 & n4249;
  assign n4251 = n805 & ~n2404;
  assign n4252 = ~n2499 & ~n4251;
  assign n4253 = n4162 & n4252;
  assign n4254 = ~n3493 & n4253;
  assign n4255 = n1278 & n4064;
  assign n4256 = n376 & n731;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~n2252 & ~n4093;
  assign n4259 = ~n3730 & n4258;
  assign n4260 = n4257 & n4259;
  assign n4261 = ~n2160 & ~n2319;
  assign n4262 = ~n2257 & n3154;
  assign n4263 = ~n891 & n4262;
  assign n4264 = n4261 & n4263;
  assign n4265 = n4260 & n4264;
  assign n4266 = n4254 & n4265;
  assign n4267 = n4250 & n4266;
  assign n4268 = ~n3068 & ~n3600;
  assign n4269 = n831 & n4268;
  assign n4270 = ~n1845 & n4269;
  assign n4271 = n3696 & n4270;
  assign n4272 = n4080 & n4271;
  assign n4273 = n4267 & n4272;
  assign n4274 = n3538 & n4273;
  assign n4275 = n2457 & n3669;
  assign po31 = ~n4274 | ~n4275;
  assign po92 = n3623 | ~n4209;
  assign n4278 = n1275 & n3495;
  assign n4279 = n4271 & n4278;
  assign po32 = po92 | ~n4279;
  assign n4281 = pi045 & pi122;
  assign n4282 = n397 & ~n4281;
  assign n4283 = ~n1464 & n3999;
  assign n4284 = n528 & n3196;
  assign n4285 = ~n4283 & ~n4284;
  assign n4286 = ~n4282 & n4285;
  assign n4287 = n3125 & n4286;
  assign n4288 = n3547 & n4287;
  assign n4289 = n974 & ~n3649;
  assign n4290 = n3648 & ~n4289;
  assign n4291 = n3785 & n4290;
  assign n4292 = pi060 & ~n379;
  assign n4293 = n381 & ~n4292;
  assign n4294 = n4223 & ~n4293;
  assign n4295 = pi014 & n2251;
  assign n4296 = ~n2288 & ~n2479;
  assign n4297 = n1262 & ~n4296;
  assign n4298 = ~n1270 & ~n4297;
  assign n4299 = ~n4295 & n4298;
  assign n4300 = n4294 & n4299;
  assign n4301 = n4291 & n4300;
  assign n4302 = n4288 & n4301;
  assign n4303 = ~pi044 & n4281;
  assign n4304 = ~n3760 & ~n4303;
  assign n4305 = n395 & ~n1914;
  assign n4306 = n236 & n4303;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = ~n4304 & ~n4307;
  assign n4309 = n4207 & ~n4308;
  assign n4310 = n3201 & n4309;
  assign n4311 = n4302 & n4310;
  assign n4312 = n4091 & n4311;
  assign n4313 = ~n1749 & ~n4024;
  assign n4314 = n3729 & n4313;
  assign n4315 = n3142 & n4314;
  assign n4316 = n2325 & n4315;
  assign n4317 = n4312 & n4316;
  assign po33 = ~n3962 | ~n4317;
  assign n4319 = n3129 & n4176;
  assign n4320 = ~n4094 & n4314;
  assign n4321 = n3752 & ~n4135;
  assign n4322 = ~n2290 & n4321;
  assign n4323 = n4320 & n4322;
  assign n4324 = ~n2668 & n4323;
  assign po34 = ~n4319 | ~n4324;
  assign n4326 = ~n287 & n2456;
  assign n4327 = n3821 & ~n4151;
  assign n4328 = n4326 & n4327;
  assign po35 = ~n3953 | ~n4328;
  assign n4330 = n4208 & n4222;
  assign n4331 = ~n938 & n4330;
  assign po36 = ~n3864 | ~n4331;
  assign n4333 = ~n2216 & ~n2317;
  assign n4334 = ~n2549 & n4333;
  assign n4335 = ~n4103 & n4334;
  assign po37 = ~n2026 | ~n4335;
  assign n4337 = ~n3494 & n3786;
  assign n4338 = n619 & ~n4113;
  assign n4339 = ~n1760 & ~n4338;
  assign n4340 = n3163 & n4339;
  assign po38 = ~n4337 | ~n4340;
  assign n4342 = n1273 & n2287;
  assign po39 = ~n2213 | ~n4342;
  assign n4344 = n2439 & n3414;
  assign n4345 = ~n2429 & ~n4344;
  assign n4346 = n540 & n4211;
  assign n4347 = n1128 & n4346;
  assign n4348 = n625 & n3848;
  assign n4349 = ~n820 & ~n4348;
  assign n4350 = ~n4347 & n4349;
  assign n4351 = ~n2688 & n4350;
  assign n4352 = ~pi045 & n2729;
  assign n4353 = ~n528 & ~n4352;
  assign n4354 = n1084 & ~n4353;
  assign n4355 = ~n1218 & ~n4354;
  assign n4356 = ~n1787 & n4355;
  assign n4357 = n4351 & n4356;
  assign n4358 = ~n1706 & ~n1760;
  assign n4359 = ~pi019 & ~n4358;
  assign n4360 = n4357 & ~n4359;
  assign n4361 = n4345 & n4360;
  assign n4362 = ~pi015 & n2237;
  assign n4363 = ~n652 & ~n4362;
  assign n4364 = ~n3545 & n4363;
  assign n4365 = ~pi039 & n1460;
  assign n4366 = n3196 & n4025;
  assign n4367 = ~n1441 & ~n4366;
  assign n4368 = ~n4365 & n4367;
  assign n4369 = ~pi044 & ~pi045;
  assign n4370 = pi122 & n4369;
  assign n4371 = n587 & n4370;
  assign n4372 = n1581 & n4371;
  assign n4373 = ~pi056 & n1213;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = ~n1975 & n4374;
  assign n4376 = n4368 & n4375;
  assign n4377 = ~n1702 & n4376;
  assign n4378 = n4364 & n4377;
  assign n4379 = n267 & n626;
  assign n4380 = ~n1664 & ~n4379;
  assign n4381 = n3827 & ~n4380;
  assign n4382 = ~pi045 & n251;
  assign n4383 = ~n385 & ~n433;
  assign n4384 = n626 & n4383;
  assign n4385 = ~n1779 & ~n4384;
  assign n4386 = ~n840 & n4385;
  assign n4387 = n4382 & ~n4386;
  assign n4388 = n1302 & n4369;
  assign n4389 = ~pi045 & n1542;
  assign n4390 = n1581 & n4389;
  assign n4391 = ~pi023 & n4382;
  assign n4392 = n373 & n4391;
  assign n4393 = ~n502 & ~n1599;
  assign n4394 = ~n1536 & n4393;
  assign n4395 = n4392 & ~n4394;
  assign n4396 = ~n4390 & ~n4395;
  assign n4397 = ~n4388 & n4396;
  assign n4398 = ~pi045 & n541;
  assign n4399 = ~n4391 & ~n4398;
  assign n4400 = n3433 & ~n4399;
  assign n4401 = n3326 & n4398;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = n4397 & n4402;
  assign n4404 = ~n4387 & n4403;
  assign n4405 = ~n4381 & n4404;
  assign n4406 = n1646 & n4398;
  assign n4407 = ~pi022 & n4382;
  assign n4408 = n662 & n4407;
  assign n4409 = ~n4406 & ~n4408;
  assign n4410 = n530 & n1170;
  assign n4411 = n4409 & ~n4410;
  assign n4412 = n382 & n1201;
  assign n4413 = ~n1197 & ~n4412;
  assign n4414 = n469 & ~n4413;
  assign n4415 = ~n2219 & ~n4414;
  assign n4416 = ~n1094 & n4415;
  assign n4417 = n4391 & ~n4416;
  assign n4418 = ~n1914 & ~n3176;
  assign n4419 = n1582 & ~n4418;
  assign n4420 = n435 & n1930;
  assign n4421 = n1445 & n4420;
  assign n4422 = ~n4419 & ~n4421;
  assign n4423 = ~n4417 & n4422;
  assign n4424 = n4411 & n4423;
  assign n4425 = ~n1930 & ~n4369;
  assign n4426 = n1305 & ~n4425;
  assign n4427 = ~n515 & n1986;
  assign n4428 = ~pi011 & n4427;
  assign n4429 = ~n4426 & ~n4428;
  assign n4430 = n3981 & n4429;
  assign n4431 = pi122 & n1579;
  assign n4432 = ~n1415 & ~n4431;
  assign n4433 = n4391 & ~n4432;
  assign n4434 = n3816 & ~n4433;
  assign n4435 = n3860 & n4434;
  assign n4436 = n4430 & n4435;
  assign n4437 = n4424 & n4436;
  assign n4438 = n4405 & n4437;
  assign n4439 = n291 & n346;
  assign n4440 = n3834 & ~n4439;
  assign n4441 = n2168 & n4440;
  assign n4442 = n977 & n3905;
  assign n4443 = n4441 & n4442;
  assign n4444 = n1059 & ~n4443;
  assign n4445 = n4438 & ~n4444;
  assign n4446 = n4378 & n4445;
  assign n4447 = n4361 & n4446;
  assign n4448 = ~pi045 & n287;
  assign n4449 = n3189 & ~n4448;
  assign n4450 = ~n3214 & n4449;
  assign n4451 = n3194 & n4179;
  assign n4452 = n4450 & n4451;
  assign n4453 = n346 & n593;
  assign n4454 = ~pi065 & n962;
  assign n4455 = ~n4453 & ~n4454;
  assign n4456 = ~n1567 & ~n1726;
  assign n4457 = ~n1413 & ~n1422;
  assign n4458 = n1564 & n4457;
  assign n4459 = n4456 & n4458;
  assign n4460 = pi122 & ~n4459;
  assign n4461 = ~n1005 & n3908;
  assign n4462 = pi065 & n855;
  assign n4463 = n1000 & n4462;
  assign n4464 = ~n1767 & ~n2662;
  assign n4465 = ~n4463 & n4464;
  assign n4466 = n4461 & n4465;
  assign n4467 = ~n4460 & n4466;
  assign n4468 = n4455 & n4467;
  assign n4469 = n956 & ~n2274;
  assign n4470 = n591 & n3884;
  assign n4471 = ~n3889 & ~n4470;
  assign n4472 = n1821 & n4471;
  assign n4473 = n290 & ~n414;
  assign n4474 = ~n628 & ~n4473;
  assign n4475 = n1618 & ~n4474;
  assign n4476 = ~n1541 & ~n4475;
  assign n4477 = n4472 & n4476;
  assign n4478 = n4469 & n4477;
  assign n4479 = n3899 & n4478;
  assign n4480 = n4468 & n4479;
  assign n4481 = ~pi045 & ~n4480;
  assign n4482 = n4452 & ~n4481;
  assign po41 = ~n4447 | ~n4482;
  assign n4484 = ~n844 & ~n3196;
  assign n4485 = n842 & ~n4484;
  assign n4486 = n1595 & n1604;
  assign n4487 = n269 & ~n4486;
  assign n4488 = ~n1366 & ~n1623;
  assign n4489 = ~n449 & ~n838;
  assign n4490 = n4488 & n4489;
  assign n4491 = ~n4487 & n4490;
  assign n4492 = ~n4485 & n4491;
  assign n4493 = n251 & n966;
  assign n4494 = n269 & n409;
  assign n4495 = ~n4493 & ~n4494;
  assign n4496 = n408 & ~n4495;
  assign n4497 = ~n389 & ~n4496;
  assign n4498 = ~pi122 & ~n3872;
  assign n4499 = ~n1245 & n1555;
  assign n4500 = ~n4498 & n4499;
  assign n4501 = ~n1639 & n4500;
  assign n4502 = ~n1576 & ~n1580;
  assign n4503 = ~n612 & n4502;
  assign n4504 = n4501 & n4503;
  assign n4505 = n4497 & n4504;
  assign n4506 = n4492 & n4505;
  assign n4507 = n3711 & n4506;
  assign n4508 = ~pi045 & ~n4507;
  assign n4509 = ~n1309 & n4369;
  assign n4510 = n343 & n3025;
  assign n4511 = n230 & n1769;
  assign n4512 = ~n3871 & ~n4511;
  assign n4513 = ~pi007 & ~n4512;
  assign n4514 = ~n4510 & ~n4513;
  assign n4515 = n1572 & n4514;
  assign n4516 = n1930 & ~n4515;
  assign n4517 = n1447 & n4420;
  assign n4518 = n773 & ~n1598;
  assign n4519 = n269 & ~n387;
  assign n4520 = ~n4518 & n4519;
  assign n4521 = ~n492 & ~n4520;
  assign n4522 = ~pi045 & n373;
  assign n4523 = ~n4521 & n4522;
  assign n4524 = ~n4517 & ~n4523;
  assign n4525 = n1548 & ~n4418;
  assign n4526 = n574 & n1769;
  assign n4527 = ~n2359 & ~n4526;
  assign n4528 = n4370 & ~n4527;
  assign n4529 = ~n4525 & ~n4528;
  assign n4530 = ~n2620 & ~n3030;
  assign n4531 = pi122 & n3848;
  assign n4532 = ~n4530 & n4531;
  assign n4533 = n1084 & n3176;
  assign n4534 = n268 & n4533;
  assign n4535 = ~n4532 & ~n4534;
  assign n4536 = n4529 & n4535;
  assign n4537 = n4524 & n4536;
  assign n4538 = n1547 & n1914;
  assign n4539 = ~n4352 & ~n4538;
  assign n4540 = n1084 & ~n4539;
  assign n4541 = pi017 & ~pi022;
  assign n4542 = n3092 & ~n4541;
  assign n4543 = n1097 & n4542;
  assign n4544 = ~n378 & ~n4543;
  assign n4545 = n4382 & ~n4544;
  assign n4546 = ~n4540 & ~n4545;
  assign n4547 = n4537 & n4546;
  assign n4548 = ~n4516 & n4547;
  assign n4549 = n4424 & n4548;
  assign n4550 = ~n4509 & n4549;
  assign n4551 = ~n4508 & n4550;
  assign n4552 = n1914 & ~n1929;
  assign n4553 = ~n3930 & n4552;
  assign n4554 = n3987 & ~n4553;
  assign n4555 = ~n1207 & n4554;
  assign n4556 = ~n575 & n3509;
  assign n4557 = ~n1233 & n4556;
  assign n4558 = ~n454 & ~n1378;
  assign n4559 = n4557 & n4558;
  assign n4560 = ~n2080 & n4559;
  assign n4561 = ~pi045 & ~n4560;
  assign n4562 = n1059 & n1935;
  assign n4563 = ~n1744 & n4562;
  assign n4564 = ~n1916 & ~n4563;
  assign n4565 = n447 & n3845;
  assign n4566 = pi021 & n4565;
  assign n4567 = ~pi056 & n1342;
  assign n4568 = n2052 & n4562;
  assign n4569 = pi004 & n4568;
  assign n4570 = ~n4567 & ~n4569;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = n528 & n2104;
  assign n4573 = n790 & n3999;
  assign n4574 = ~pi061 & pi065;
  assign n4575 = n534 & n4574;
  assign n4576 = n1312 & n4575;
  assign n4577 = n284 & n4576;
  assign n4578 = ~n4573 & ~n4577;
  assign n4579 = ~n4572 & n4578;
  assign n4580 = ~n4008 & n4579;
  assign n4581 = n4571 & n4580;
  assign n4582 = n4564 & n4581;
  assign n4583 = n4285 & n4582;
  assign n4584 = ~n4561 & n4583;
  assign n4585 = n4555 & n4584;
  assign n4586 = n502 & n2584;
  assign n4587 = n386 & n662;
  assign n4588 = ~n775 & ~n4587;
  assign n4589 = ~n4586 & n4588;
  assign n4590 = ~n2581 & n4589;
  assign n4591 = ~n725 & ~n856;
  assign n4592 = n376 & ~n4591;
  assign n4593 = n774 & n2517;
  assign n4594 = ~n1408 & n2572;
  assign n4595 = n1126 & n4594;
  assign n4596 = ~n2538 & ~n4595;
  assign n4597 = ~n4593 & n4596;
  assign n4598 = ~n4592 & n4597;
  assign n4599 = n4590 & n4598;
  assign n4600 = n2965 & n4599;
  assign n4601 = n2566 & n4600;
  assign n4602 = n1132 & n3900;
  assign n4603 = ~n1767 & n4602;
  assign n4604 = ~pi045 & ~n4603;
  assign n4605 = ~pi045 & n3913;
  assign n4606 = n774 & n4392;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4604 & n4607;
  assign n4609 = n735 & n855;
  assign n4610 = n672 & n4346;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n2897 & n4611;
  assign n4613 = ~pi023 & n735;
  assign n4614 = ~n731 & ~n4613;
  assign n4615 = n1197 & ~n4614;
  assign n4616 = n518 & n3983;
  assign n4617 = ~n1089 & n4616;
  assign n4618 = ~pi122 & n1154;
  assign n4619 = ~n1415 & ~n1942;
  assign n4620 = ~n4618 & n4619;
  assign n4621 = n4391 & ~n4620;
  assign n4622 = ~n1877 & ~n3979;
  assign n4623 = ~n4621 & n4622;
  assign n4624 = ~n4617 & n4623;
  assign n4625 = ~n4615 & n4624;
  assign n4626 = n4612 & n4625;
  assign n4627 = n4608 & n4626;
  assign n4628 = n4601 & n4627;
  assign n4629 = ~n1154 & ~n2742;
  assign n4630 = n251 & ~n4629;
  assign n4631 = n1418 & ~n1745;
  assign n4632 = n1921 & n4631;
  assign n4633 = n4457 & n4632;
  assign n4634 = ~n4630 & n4633;
  assign n4635 = n1930 & ~n4634;
  assign n4636 = n268 & n3903;
  assign n4637 = n1930 & n4636;
  assign n4638 = ~n2563 & ~n4637;
  assign n4639 = n1151 & n4346;
  assign n4640 = ~pi122 & n4639;
  assign n4641 = n1428 & n2358;
  assign n4642 = ~pi045 & n4641;
  assign n4643 = ~pi003 & n4642;
  assign n4644 = n269 & n1848;
  assign n4645 = n346 & n3840;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~n4643 & n4646;
  assign n4648 = ~n738 & ~n1536;
  assign n4649 = ~n569 & n4648;
  assign n4650 = n1217 & ~n4649;
  assign n4651 = n4647 & ~n4650;
  assign n4652 = ~n4640 & n4651;
  assign n4653 = ~pi021 & n2560;
  assign n4654 = n452 & n4653;
  assign n4655 = ~n2696 & ~n4654;
  assign n4656 = ~n4427 & n4655;
  assign n4657 = n4652 & n4656;
  assign n4658 = n4638 & n4657;
  assign n4659 = ~n631 & n4658;
  assign n4660 = ~n4635 & n4659;
  assign n4661 = n4378 & n4660;
  assign n4662 = n4628 & n4661;
  assign n4663 = ~n396 & ~n4052;
  assign n4664 = ~po67 & n2264;
  assign n4665 = n1455 & n4664;
  assign n4666 = n4663 & n4665;
  assign n4667 = ~n608 & n1145;
  assign n4668 = ~n1726 & n3915;
  assign n4669 = n4667 & n4668;
  assign n4670 = n4666 & n4669;
  assign n4671 = ~n2055 & n4670;
  assign n4672 = n3909 & n4469;
  assign n4673 = n4671 & n4672;
  assign n4674 = ~pi045 & ~n4673;
  assign n4675 = n4662 & ~n4674;
  assign n4676 = n4585 & n4675;
  assign n4677 = n4551 & n4676;
  assign n4678 = n3865 & n4677;
  assign n4679 = ~n3784 & n4358;
  assign n4680 = ~pi011 & n2161;
  assign n4681 = n2442 & ~n4680;
  assign n4682 = pi065 & n2423;
  assign n4683 = ~n2422 & ~n4682;
  assign n4684 = ~n3238 & n4683;
  assign n4685 = n4681 & n4684;
  assign n4686 = n4679 & n4685;
  assign n4687 = pi012 & ~n4247;
  assign n4688 = ~n2446 & ~n4687;
  assign n4689 = ~n654 & n2886;
  assign n4690 = ~n3386 & ~n4689;
  assign n4691 = n2484 & n4690;
  assign n4692 = n4688 & n4691;
  assign n4693 = pi012 & n911;
  assign n4694 = n3533 & ~n4693;
  assign n4695 = ~n3152 & n3341;
  assign n4696 = n866 & ~n4695;
  assign n4697 = pi023 & ~n2455;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = n4694 & n4698;
  assign n4700 = n2495 & ~n2612;
  assign n4701 = ~n713 & n4700;
  assign n4702 = ~n2336 & n4701;
  assign n4703 = n4699 & n4702;
  assign n4704 = n2451 & n4703;
  assign n4705 = ~n4093 & n4704;
  assign n4706 = n4692 & n4705;
  assign n4707 = n4686 & n4706;
  assign n4708 = n1305 & n3176;
  assign n4709 = n1046 & n1059;
  assign n4710 = n3176 & n3888;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = ~n4708 & n4711;
  assign n4713 = n702 & n1748;
  assign n4714 = ~n4115 & n4148;
  assign n4715 = n1059 & ~n4714;
  assign n4716 = n1914 & n3904;
  assign n4717 = ~n4715 & ~n4716;
  assign n4718 = ~n4713 & n4717;
  assign n4719 = n3995 & n4718;
  assign n4720 = n1789 & n4719;
  assign n4721 = n4712 & n4720;
  assign n4722 = n4707 & n4721;
  assign n4723 = n922 & n4129;
  assign n4724 = ~n4134 & ~n4723;
  assign n4725 = n4113 & ~n4724;
  assign n4726 = n283 & n4123;
  assign n4727 = ~n284 & ~n4726;
  assign n4728 = ~n4725 & ~n4727;
  assign n4729 = n619 & n4124;
  assign n4730 = n584 & n766;
  assign n4731 = n4125 & ~n4730;
  assign n4732 = ~n922 & n4132;
  assign n4733 = n4130 & ~n4732;
  assign n4734 = ~n336 & ~n1085;
  assign n4735 = n4117 & n4734;
  assign n4736 = ~n4733 & ~n4735;
  assign n4737 = ~n4731 & n4736;
  assign n4738 = n1059 & ~n4737;
  assign n4739 = ~n4729 & ~n4738;
  assign n4740 = ~n4728 & n4739;
  assign n4741 = n4722 & n4740;
  assign po42 = ~n4678 | ~n4741;
  assign n4743 = ~n411 & n1269;
  assign n4744 = n343 & ~n4743;
  assign n4745 = n2054 & ~n4744;
  assign n4746 = ~n573 & ~n1470;
  assign n4747 = ~n1800 & n4746;
  assign n4748 = n343 & ~n4747;
  assign n4749 = n372 & n1065;
  assign n4750 = ~n638 & ~n1312;
  assign n4751 = ~n4749 & n4750;
  assign n4752 = ~n4748 & n4751;
  assign n4753 = n4714 & n4752;
  assign n4754 = n992 & n4753;
  assign n4755 = n4745 & n4754;
  assign n4756 = n1059 & ~n4755;
  assign n4757 = ~pi006 & n4637;
  assign n4758 = n2371 & n3856;
  assign n4759 = n1044 & n4758;
  assign n4760 = ~n4642 & ~n4759;
  assign n4761 = ~n3238 & ~n4217;
  assign n4762 = n4760 & n4761;
  assign n4763 = ~n4757 & n4762;
  assign n4764 = n1028 & ~n4418;
  assign n4765 = ~n4710 & ~n4764;
  assign n4766 = n4763 & n4765;
  assign n4767 = n949 & n4392;
  assign n4768 = n4537 & ~n4767;
  assign n4769 = ~n2438 & n4768;
  assign n4770 = ~n1631 & n1666;
  assign n4771 = ~n1385 & n4770;
  assign n4772 = n3827 & ~n4771;
  assign n4773 = n4769 & ~n4772;
  assign n4774 = n3820 & n4773;
  assign n4775 = n3852 & n4774;
  assign n4776 = n4766 & n4775;
  assign n4777 = n4585 & n4776;
  assign n4778 = n4345 & n4740;
  assign n4779 = n4777 & n4778;
  assign n4780 = ~n4756 & n4779;
  assign n4781 = n1029 & n3175;
  assign n4782 = n1047 & n4369;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = ~n3992 & n4783;
  assign n4785 = n4450 & n4784;
  assign n4786 = n4492 & n4666;
  assign n4787 = pi065 & n962;
  assign n4788 = ~n753 & n1639;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = n1000 & n1001;
  assign n4791 = n411 & n540;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = n4789 & n4792;
  assign n4794 = n609 & n2303;
  assign n4795 = ~n4494 & ~n4794;
  assign n4796 = ~n1136 & n4795;
  assign n4797 = n408 & ~n4796;
  assign n4798 = ~n3914 & ~n4797;
  assign n4799 = ~n1673 & n4798;
  assign n4800 = ~n591 & n3883;
  assign n4801 = ~n2358 & ~n4800;
  assign n4802 = n560 & ~n4801;
  assign n4803 = ~n2408 & ~n4802;
  assign n4804 = ~n571 & n4803;
  assign n4805 = ~n1637 & n4804;
  assign n4806 = ~pi044 & ~n4225;
  assign n4807 = ~pi122 & n4526;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = n1555 & n4808;
  assign n4810 = n4805 & n4809;
  assign n4811 = n4799 & n4810;
  assign n4812 = n3824 & n4811;
  assign n4813 = n4793 & n4812;
  assign n4814 = n4786 & n4813;
  assign n4815 = ~pi045 & ~n4814;
  assign n4816 = n540 & n1154;
  assign n4817 = n1570 & n4632;
  assign n4818 = ~n4816 & n4817;
  assign n4819 = n1930 & ~n4818;
  assign n4820 = ~n4815 & ~n4819;
  assign n4821 = n4785 & n4820;
  assign po43 = ~n4780 | ~n4821;
  assign n4823 = ~n3525 & ~n4241;
  assign n4824 = n394 & n1152;
  assign n4825 = ~n2561 & ~n4824;
  assign n4826 = n4601 & n4825;
  assign n4827 = n4823 & n4826;
  assign po44 = ~n4707 | ~n4827;
  assign po45 = ~n4452 | ~n4686;
  assign n4830 = n4685 & n4785;
  assign n4831 = ~n4177 & n4765;
  assign n4832 = ~n3193 & n4831;
  assign n4833 = ~n1749 & ~n4716;
  assign n4834 = ~n4708 & n4833;
  assign n4835 = ~n1787 & n4834;
  assign n4836 = n4832 & n4835;
  assign n4837 = n4830 & n4836;
  assign po46 = ~n4678 | ~n4837;
  assign n4839 = n284 & ~n4113;
  assign n4840 = ~n1787 & ~n4839;
  assign n4841 = ~n2697 & n4840;
  assign po47 = ~n4679 | ~n4841;
  assign n4843 = pi004 & n2025;
  assign n4844 = ~n3546 & ~n4843;
  assign po49 = ~n4368 | n4844;
  assign n4846 = n284 & n4724;
  assign n4847 = ~n1702 & ~n4846;
  assign po50 = ~n4681 | ~n4847;
  assign n4849 = pi026 & n4726;
  assign n4850 = ~n4729 & ~n4849;
  assign n4851 = ~n1975 & n4850;
  assign po51 = ~n4622 | ~n4851;
  assign n4853 = ~n2462 & n2631;
  assign n4854 = ~n874 & n4853;
  assign po52 = n4693 | ~n4854;
  assign n4856 = ~n2882 & n4692;
  assign po53 = n2635 | ~n4856;
  assign n4858 = ~n4373 & ~n4567;
  assign n4859 = ~n2336 & n4858;
  assign n4860 = ~n2353 & ~n4410;
  assign n4861 = n4859 & n4860;
  assign po54 = ~n3821 | ~n4861;
  assign n4863 = n1155 & ~n1415;
  assign n4864 = n4391 & ~n4863;
  assign n4865 = pi039 & pi045;
  assign n4866 = ~pi122 & n4865;
  assign n4867 = n343 & n1063;
  assign n4868 = n632 & n1096;
  assign n4869 = ~n4867 & ~n4868;
  assign n4870 = ~n2407 & n4869;
  assign n4871 = n4866 & ~n4870;
  assign n4872 = ~n4639 & ~n4871;
  assign n4873 = n1214 & n4872;
  assign n4874 = n235 & n3999;
  assign n4875 = ~n4610 & ~n4874;
  assign n4876 = n4712 & n4875;
  assign n4877 = n4873 & n4876;
  assign n4878 = ~n395 & n4669;
  assign n4879 = ~n454 & n4878;
  assign n4880 = n3910 & n4879;
  assign n4881 = ~pi045 & ~n4880;
  assign n4882 = n4551 & ~n4881;
  assign n4883 = n4877 & n4882;
  assign n4884 = n4608 & n4883;
  assign n4885 = ~n4864 & n4884;
  assign n4886 = ~n3176 & ~n3938;
  assign n4887 = n3171 & ~n4886;
  assign n4888 = n3948 & ~n4887;
  assign n4889 = ~n3937 & n4886;
  assign n4890 = ~n1033 & ~n4889;
  assign n4891 = n311 & ~n1029;
  assign n4892 = ~n355 & n4891;
  assign n4893 = ~n3941 & ~n4892;
  assign n4894 = ~n3170 & ~n3940;
  assign n4895 = ~n4893 & ~n4894;
  assign n4896 = ~n4890 & n4895;
  assign n4897 = n4888 & n4896;
  assign n4898 = ~n1032 & ~n3941;
  assign n4899 = ~n3951 & ~n4898;
  assign n4900 = n4897 & n4899;
  assign n4901 = ~n4372 & ~n4566;
  assign n4902 = ~n2500 & n4901;
  assign n4903 = n375 & n4565;
  assign n4904 = n4902 & ~n4903;
  assign n4905 = n4900 & n4904;
  assign po57 = ~n4885 | ~n4905;
  assign n4907 = ~n2910 & ~n4427;
  assign n4908 = ~pi011 & ~n4907;
  assign po55 = po57 | n4908;
  assign n4910 = pi020 & po67;
  assign n4911 = n2421 & n4462;
  assign n4912 = ~pi018 & ~n729;
  assign n4913 = n394 & ~n4912;
  assign n4914 = ~n409 & n4913;
  assign n4915 = n230 & n2303;
  assign n4916 = ~n4073 & ~n4915;
  assign n4917 = ~n386 & n4916;
  assign n4918 = ~n4914 & n4917;
  assign n4919 = n277 & ~n4918;
  assign n4920 = ~n4911 & ~n4919;
  assign n4921 = ~n4910 & n4920;
  assign n4922 = n714 & n4921;
  assign po58 = n938 | ~n4922;
  assign po56 = ~n4907 | po58;
  assign po59 = po57 | n4911;
  assign n4926 = ~pi020 & n1643;
  assign n4927 = ~n3433 & ~n4926;
  assign n4928 = n609 & ~n4927;
  assign n4929 = ~pi044 & n393;
  assign n4930 = ~n643 & ~n4929;
  assign n4931 = ~n1825 & n4930;
  assign n4932 = n541 & ~n4931;
  assign n4933 = ~n4928 & ~n4932;
  assign n4934 = n1930 & ~n4933;
  assign n4935 = n542 & n3344;
  assign n4936 = ~n3678 & ~n4935;
  assign n4937 = n3176 & ~n4936;
  assign n4938 = ~n382 & n4606;
  assign n4939 = ~n4371 & ~n4389;
  assign n4940 = n1283 & ~n4939;
  assign n4941 = ~n4938 & ~n4940;
  assign n4942 = ~n4621 & n4941;
  assign n4943 = ~n4937 & n4942;
  assign n4944 = pi122 & ~n1651;
  assign n4945 = ~n1131 & n4944;
  assign n4946 = n4604 & ~n4945;
  assign n4947 = n3911 & n4391;
  assign n4948 = n4907 & ~n4947;
  assign n4949 = n4920 & n4948;
  assign n4950 = ~n4946 & n4949;
  assign n4951 = n4943 & n4950;
  assign n4952 = ~n4934 & n4951;
  assign n4953 = n4883 & n4952;
  assign po60 = ~n4905 | ~n4953;
  assign n4955 = ~n4410 & n4900;
  assign po61 = n1213 | ~n4955;
  assign n4957 = ~n2751 & n3046;
  assign n4958 = n2234 & n4957;
  assign n4959 = ~n2181 & ~n2544;
  assign n4960 = pi013 & n1158;
  assign n4961 = ~n2131 & ~n4960;
  assign n4962 = ~n2680 & n4961;
  assign n4963 = n4959 & n4962;
  assign n4964 = n3563 & n4963;
  assign po62 = ~n4958 | ~n4964;
  assign n4966 = n398 & ~n1250;
  assign n4967 = n973 & ~n1070;
  assign n4968 = n969 & ~n1070;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = ~n266 & n4969;
  assign n4971 = ~n990 & ~n1070;
  assign n4972 = n4970 & ~n4971;
  assign n4973 = ~n1075 & ~n1348;
  assign n4974 = ~n1521 & ~n3082;
  assign n4975 = n4973 & n4974;
  assign n4976 = ~n3511 & n4975;
  assign n4977 = ~n635 & n4976;
  assign n4978 = n371 & ~n1070;
  assign n4979 = ~n3277 & ~n4978;
  assign n4980 = n1331 & n1469;
  assign n4981 = n4979 & ~n4980;
  assign n4982 = n1025 & n4981;
  assign n4983 = n1435 & n4982;
  assign n4984 = n4977 & n4983;
  assign n4985 = n4972 & n4984;
  assign n4986 = n4966 & n4985;
  assign n4987 = n301 & ~n1039;
  assign n4988 = n2158 & n4987;
  assign n4989 = n606 & n4988;
  assign po63 = ~n4986 | ~n4989;
  assign n4991 = ~n1943 & n2946;
  assign n4992 = pi019 & n2927;
  assign n4993 = ~n1092 & ~n4992;
  assign n4994 = n2916 & n4993;
  assign n4995 = ~n1697 & n4994;
  assign n4996 = ~n1656 & n4995;
  assign n4997 = n1560 & n4996;
  assign n4998 = n1294 & n2679;
  assign po65 = n3554 | ~n4998;
  assign n5000 = ~pi039 & n4517;
  assign n5001 = n3086 & ~n5000;
  assign n5002 = ~n1612 & ~n2903;
  assign n5003 = ~n1467 & n5002;
  assign n5004 = n2684 & n5003;
  assign n5005 = n757 & n1215;
  assign n5006 = n5004 & n5005;
  assign n5007 = n5001 & n5006;
  assign n5008 = ~po65 & n5007;
  assign n5009 = n4997 & n5008;
  assign n5010 = n4991 & n5009;
  assign n5011 = n2221 & n5010;
  assign n5012 = ~n1366 & ~n2894;
  assign n5013 = n1485 & n5012;
  assign n5014 = n1289 & n5013;
  assign n5015 = ~n383 & n1229;
  assign n5016 = ~n1446 & ~n5015;
  assign n5017 = n5014 & n5016;
  assign n5018 = n3067 & n5017;
  assign n5019 = n1058 & n5018;
  assign po64 = ~n5011 | ~n5019;
  assign po66 = n938 | ~n3743;
  assign n5022 = pi013 & n1905;
  assign n5023 = ~n356 & ~n5022;
  assign n5024 = ~n1976 & n5023;
  assign n5025 = ~n1023 & ~n2777;
  assign n5026 = ~n3222 & n5025;
  assign po68 = ~n5024 | ~n5026;
  assign n5028 = pi065 & n2419;
  assign n5029 = ~pi010 & n2446;
  assign n5030 = ~n1760 & ~n5029;
  assign n5031 = ~n5028 & n5030;
  assign n5032 = ~n2422 & ~po48;
  assign n5033 = ~n1611 & n5032;
  assign n5034 = n5024 & n5033;
  assign n5035 = ~pi023 & n2454;
  assign n5036 = ~pi018 & n2459;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = n1024 & n4854;
  assign n5039 = n5037 & n5038;
  assign n5040 = n5034 & n5039;
  assign n5041 = n5031 & n5040;
  assign n5042 = n1308 & n3743;
  assign n5043 = n1237 & ~n2500;
  assign n5044 = n5042 & n5043;
  assign n5045 = n1598 & n1607;
  assign n5046 = ~n3784 & ~n5045;
  assign n5047 = pi012 & ~n919;
  assign n5048 = n2478 & ~n5047;
  assign n5049 = n5046 & n5048;
  assign n5050 = n5044 & n5049;
  assign po69 = ~n5041 | ~n5050;
  assign po70 = n3481 | n5028;
  assign n5053 = n337 & n3903;
  assign n5054 = pi004 & n2316;
  assign n5055 = ~n5053 & ~n5054;
  assign n5056 = ~n2139 & n5055;
  assign n5057 = ~n2146 & ~n2312;
  assign n5058 = ~n2004 & n5057;
  assign n5059 = n5056 & n5058;
  assign n5060 = pi108 & ~n5059;
  assign n5061 = ~n1178 & ~n5060;
  assign n5062 = pi061 & pi122;
  assign n5063 = ~pi062 & ~n5062;
  assign n5064 = n551 & n3196;
  assign n5065 = ~n1159 & ~n5064;
  assign n5066 = ~pi031 & ~n5065;
  assign n5067 = ~n5063 & n5066;
  assign n5068 = ~n1380 & ~n4365;
  assign n5069 = ~pi031 & ~n5068;
  assign n5070 = ~pi032 & n5069;
  assign n5071 = ~n5067 & ~n5070;
  assign n5072 = pi039 & n2095;
  assign n5073 = pi033 & n5072;
  assign n5074 = n1019 & ~n2129;
  assign n5075 = ~n5073 & n5074;
  assign n5076 = pi060 & n1061;
  assign n5077 = ~n1509 & ~n5076;
  assign n5078 = n5075 & n5077;
  assign n5079 = n300 & n5078;
  assign n5080 = ~n3558 & n5079;
  assign n5081 = n5071 & n5080;
  assign n5082 = n5061 & n5081;
  assign n5083 = ~pi039 & ~n4564;
  assign n5084 = ~pi045 & n2215;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = pi061 & ~pi062;
  assign n5087 = pi039 & n3275;
  assign n5088 = ~pi031 & n5087;
  assign n5089 = ~n5086 & n5088;
  assign n5090 = ~n887 & ~n5089;
  assign n5091 = n5085 & n5090;
  assign n5092 = n5082 & n5091;
  assign n5093 = ~n1920 & ~n3927;
  assign n5094 = n1930 & ~n5093;
  assign n5095 = n5092 & ~n5094;
  assign n5096 = pi097 & ~n1506;
  assign n5097 = pi031 & pi039;
  assign n5098 = n1460 & n5097;
  assign n5099 = ~n2191 & ~n5098;
  assign n5100 = ~n617 & n5099;
  assign n5101 = n1922 & n1935;
  assign n5102 = pi051 & n5101;
  assign n5103 = n5100 & ~n5102;
  assign n5104 = ~n5096 & n5103;
  assign n5105 = n539 & ~n2011;
  assign n5106 = ~n2422 & n5105;
  assign n5107 = n1920 & n1935;
  assign n5108 = n1918 & ~n3931;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = pi045 & ~n5109;
  assign n5111 = ~n2262 & ~n5072;
  assign n5112 = ~n688 & n5111;
  assign n5113 = pi034 & ~n5112;
  assign n5114 = ~n5110 & ~n5113;
  assign n5115 = n5106 & n5114;
  assign n5116 = ~n4968 & n5115;
  assign n5117 = ~n957 & n5116;
  assign n5118 = ~n1314 & ~n1348;
  assign n5119 = ~n2419 & n5118;
  assign n5120 = ~n427 & n5119;
  assign n5121 = ~n3081 & n5120;
  assign n5122 = pi065 & ~n5121;
  assign n5123 = n692 & n2082;
  assign n5124 = pi092 & n879;
  assign n5125 = n1501 & n5124;
  assign n5126 = ~n5123 & ~n5125;
  assign n5127 = pi109 & n4035;
  assign n5128 = ~n2149 & ~n2316;
  assign n5129 = n5127 & ~n5128;
  assign n5130 = n1915 & n1920;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = n5126 & n5131;
  assign n5133 = ~n5122 & n5132;
  assign n5134 = n2451 & n5133;
  assign n5135 = ~n1937 & n4865;
  assign n5136 = ~pi045 & n3932;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = ~n3931 & ~n5137;
  assign n5139 = n5134 & ~n5138;
  assign n5140 = n5117 & n5139;
  assign n5141 = n5104 & n5140;
  assign po71 = ~n5095 | ~n5141;
  assign n5143 = n1109 & n2596;
  assign n5144 = n369 & n4653;
  assign n5145 = ~n5143 & ~n5144;
  assign n5146 = n4590 & n5145;
  assign n5147 = ~n2518 & n5146;
  assign n5148 = pi076 & ~n5147;
  assign n5149 = ~pi077 & ~n745;
  assign n5150 = ~n249 & ~n321;
  assign n5151 = ~n302 & ~n5150;
  assign n5152 = ~pi058 & ~pi059;
  assign n5153 = n2307 & ~n5152;
  assign n5154 = ~n5151 & ~n5153;
  assign n5155 = ~n5149 & n5154;
  assign n5156 = ~pi040 & ~pi041;
  assign n5157 = ~n2247 & ~n5156;
  assign n5158 = n3705 & ~n5157;
  assign n5159 = n284 & n2050;
  assign n5160 = ~pi032 & pi039;
  assign n5161 = n1460 & n5160;
  assign n5162 = ~n5159 & ~n5161;
  assign n5163 = ~n2117 & n5162;
  assign n5164 = ~pi031 & ~n5163;
  assign n5165 = n1931 & ~n3933;
  assign n5166 = n2015 & ~n5165;
  assign n5167 = ~n5164 & n5166;
  assign n5168 = n5158 & n5167;
  assign n5169 = n5155 & n5168;
  assign n5170 = ~n5148 & n5169;
  assign n5171 = n1928 & ~n1936;
  assign n5172 = ~n1747 & ~n5171;
  assign n5173 = ~pi039 & ~n5172;
  assign n5174 = ~n1918 & ~n1923;
  assign n5175 = ~n1401 & n5174;
  assign n5176 = ~n1926 & ~n5175;
  assign n5177 = n2151 & ~n3929;
  assign n5178 = ~n5176 & n5177;
  assign n5179 = ~n5173 & n5178;
  assign n5180 = ~n383 & n4463;
  assign n5181 = n1220 & ~n5180;
  assign n5182 = n5179 & n5181;
  assign n5183 = n5170 & n5182;
  assign n5184 = ~n4004 & ~n5097;
  assign n5185 = n572 & ~n5184;
  assign n5186 = ~pi052 & n2567;
  assign n5187 = pi049 & n5186;
  assign n5188 = ~n5185 & ~n5187;
  assign n5189 = ~n2129 & ~n2309;
  assign n5190 = ~n2650 & n5189;
  assign n5191 = pi108 & ~n5190;
  assign n5192 = ~n4967 & ~n5191;
  assign n5193 = n5188 & n5192;
  assign n5194 = pi051 & pi089;
  assign n5195 = n2669 & n5194;
  assign n5196 = pi065 & n3019;
  assign n5197 = ~n3277 & ~n5196;
  assign n5198 = ~n2452 & ~n2812;
  assign n5199 = n5197 & n5198;
  assign n5200 = ~n5195 & n5199;
  assign n5201 = ~n619 & n1070;
  assign n5202 = n2449 & ~n5201;
  assign n5203 = n5200 & ~n5202;
  assign n5204 = n5193 & n5203;
  assign n5205 = ~pi051 & pi089;
  assign n5206 = n2461 & ~n5205;
  assign n5207 = n892 & n5206;
  assign n5208 = ~pi051 & pi088;
  assign n5209 = ~n1849 & ~n5208;
  assign n5210 = pi006 & n5209;
  assign n5211 = n2093 & n5210;
  assign n5212 = ~n5107 & ~n5211;
  assign n5213 = ~n5207 & n5212;
  assign n5214 = pi061 & ~pi122;
  assign n5215 = ~n591 & n5214;
  assign n5216 = ~pi005 & n5215;
  assign n5217 = ~n223 & n5062;
  assign n5218 = n345 & n5217;
  assign n5219 = ~n5216 & ~n5218;
  assign n5220 = n426 & ~n5219;
  assign n5221 = ~n2654 & ~n5220;
  assign n5222 = pi074 & n1757;
  assign n5223 = pi050 & ~pi051;
  assign n5224 = n2917 & ~n5223;
  assign n5225 = ~n1896 & ~n5224;
  assign n5226 = ~n5222 & n5225;
  assign n5227 = n5221 & n5226;
  assign n5228 = ~pi034 & n5073;
  assign n5229 = ~pi106 & n1390;
  assign n5230 = pi048 & ~pi051;
  assign n5231 = ~pi077 & n5230;
  assign n5232 = ~pi014 & n2029;
  assign n5233 = ~n5231 & n5232;
  assign n5234 = ~n5229 & ~n5233;
  assign n5235 = ~n5228 & n5234;
  assign n5236 = pi104 & n1378;
  assign n5237 = ~n3091 & ~n5236;
  assign n5238 = n5235 & n5237;
  assign n5239 = n2721 & n5238;
  assign n5240 = n5227 & n5239;
  assign n5241 = n5213 & n5240;
  assign n5242 = n5204 & n5241;
  assign n5243 = ~pi062 & ~n5214;
  assign n5244 = n5088 & ~n5243;
  assign n5245 = n5104 & ~n5244;
  assign n5246 = n5242 & n5245;
  assign n5247 = n5183 & n5246;
  assign n5248 = ~pi066 & ~n4843;
  assign n5249 = ~n2026 & n5248;
  assign n5250 = ~n2589 & ~n5249;
  assign n5251 = n336 & n5127;
  assign n5252 = n269 & ~n1935;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = n3903 & ~n5253;
  assign n5255 = n695 & n2082;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = pi105 & n481;
  assign n5258 = ~n2027 & ~n5257;
  assign n5259 = ~n1518 & n5258;
  assign n5260 = n5256 & n5259;
  assign n5261 = ~n1617 & n5260;
  assign n5262 = ~pi090 & n1501;
  assign n5263 = pi091 & n5262;
  assign n5264 = ~n3803 & ~n5263;
  assign n5265 = n1511 & n5264;
  assign n5266 = n5261 & n5265;
  assign n5267 = pi027 & n2449;
  assign n5268 = pi045 & n2068;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = n282 & ~n5269;
  assign n5271 = n5266 & ~n5270;
  assign n5272 = n5250 & n5271;
  assign n5273 = pi032 & n5069;
  assign n5274 = pi067 & ~n3959;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = n5066 & n5243;
  assign n5277 = pi034 & n692;
  assign n5278 = pi027 & n302;
  assign n5279 = ~pi108 & n353;
  assign n5280 = ~n5278 & n5279;
  assign n5281 = ~n350 & n5280;
  assign n5282 = ~n5277 & ~n5281;
  assign n5283 = ~n4911 & n5282;
  assign n5284 = ~n5276 & n5283;
  assign n5285 = ~n4682 & n5284;
  assign n5286 = n5275 & n5285;
  assign n5287 = n5272 & n5286;
  assign n5288 = n1315 & n1342;
  assign n5289 = n5119 & ~n5288;
  assign n5290 = ~n639 & ~n1340;
  assign n5291 = n5289 & n5290;
  assign n5292 = ~n1471 & n5291;
  assign n5293 = pi061 & ~n5292;
  assign n5294 = n3991 & ~n5293;
  assign n5295 = n5287 & n5294;
  assign po72 = ~n5247 | ~n5295;
  assign n5297 = ~n1061 & ~n1617;
  assign n5298 = ~n3021 & n4979;
  assign n5299 = n3661 & n5298;
  assign po73 = ~n5297 | ~n5299;
  assign n5301 = ~n401 & ~n3762;
  assign n5302 = ~n1437 & n5301;
  assign n5303 = n5299 & n5302;
  assign n5304 = n947 & n1545;
  assign n5305 = pi021 & n5304;
  assign n5306 = ~n1638 & ~n5305;
  assign n5307 = n5303 & n5306;
  assign n5308 = ~n526 & n620;
  assign n5309 = ~n1070 & n4749;
  assign n5310 = ~n3601 & ~n5309;
  assign n5311 = n5297 & n5310;
  assign n5312 = ~n5308 & n5311;
  assign n5313 = n1081 & n5312;
  assign po77 = ~n5307 | ~n5313;
  assign n5315 = n588 & n643;
  assign n5316 = n472 & n672;
  assign n5317 = ~n1525 & ~n5316;
  assign n5318 = ~n410 & n5317;
  assign n5319 = ~n3437 & n5318;
  assign n5320 = n843 & ~n5319;
  assign n5321 = ~n1282 & ~n4226;
  assign n5322 = ~n2695 & n5321;
  assign n5323 = n1183 & n1187;
  assign n5324 = ~n465 & ~n1119;
  assign n5325 = ~n5323 & n5324;
  assign n5326 = pi023 & n1536;
  assign n5327 = n1607 & ~n5326;
  assign n5328 = pi019 & n5327;
  assign n5329 = ~n1387 & ~n5328;
  assign n5330 = n5325 & n5329;
  assign n5331 = n5322 & n5330;
  assign n5332 = ~n5320 & n5331;
  assign n5333 = ~n5315 & n5332;
  assign n5334 = pi003 & n2357;
  assign n5335 = ~n2363 & ~n5334;
  assign n5336 = ~n1546 & n2753;
  assign n5337 = ~n5335 & n5336;
  assign n5338 = ~n1286 & n5337;
  assign n5339 = ~n1101 & n1624;
  assign n5340 = ~n614 & n5339;
  assign n5341 = n5338 & n5340;
  assign n5342 = ~n372 & ~n1109;
  assign n5343 = n1806 & ~n5342;
  assign n5344 = n5341 & ~n5343;
  assign n5345 = n5333 & n5344;
  assign n5346 = ~po00 & n5303;
  assign n5347 = n1077 & ~n2909;
  assign n5348 = ~n1078 & n5347;
  assign n5349 = n5346 & n5348;
  assign n5350 = n457 & ~n504;
  assign n5351 = ~pi019 & ~n5350;
  assign n5352 = n748 & n1193;
  assign n5353 = ~n383 & n5352;
  assign n5354 = ~n5351 & ~n5353;
  assign n5355 = n5349 & n5354;
  assign n5356 = n2789 & n5355;
  assign po78 = ~n5345 | ~n5356;
  assign n5358 = ~n1386 & ~n1476;
  assign n5359 = n505 & n5358;
  assign n5360 = n3576 & n5359;
  assign n5361 = ~pi122 & n1083;
  assign n5362 = n1553 & ~n5361;
  assign n5363 = ~n3914 & ~n5362;
  assign n5364 = ~n1138 & n3891;
  assign n5365 = n3432 & n5364;
  assign n5366 = n5363 & n5365;
  assign n5367 = ~n383 & ~n5366;
  assign n5368 = n5346 & ~n5367;
  assign n5369 = n5360 & n5368;
  assign n5370 = n1809 & n3042;
  assign n5371 = ~n2780 & n5370;
  assign n5372 = n5338 & n5371;
  assign n5373 = n5369 & n5372;
  assign n5374 = ~n1675 & n3244;
  assign n5375 = n588 & ~n5374;
  assign n5376 = ~n1964 & ~n5375;
  assign n5377 = n1089 & n1481;
  assign n5378 = ~n1283 & ~n1581;
  assign n5379 = ~n3673 & ~n5378;
  assign n5380 = ~n5377 & ~n5379;
  assign n5381 = n5376 & n5380;
  assign n5382 = ~n1536 & ~n2850;
  assign n5383 = n1281 & ~n5382;
  assign n5384 = ~n1648 & ~n5383;
  assign n5385 = n2202 & n5384;
  assign n5386 = n3215 & n5385;
  assign n5387 = n583 & n800;
  assign n5388 = ~pi020 & n3059;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = ~n1302 & n5389;
  assign n5391 = n1615 & n5390;
  assign n5392 = n5386 & n5391;
  assign n5393 = n224 & n392;
  assign n5394 = ~pi122 & n373;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = n492 & ~n5395;
  assign n5397 = ~pi018 & n1862;
  assign n5398 = ~n277 & ~n471;
  assign n5399 = ~n1778 & n5398;
  assign n5400 = n5397 & ~n5399;
  assign n5401 = ~n5396 & ~n5400;
  assign n5402 = pi003 & n1551;
  assign n5403 = ~n1638 & ~n5402;
  assign n5404 = n5401 & n5403;
  assign n5405 = ~n1242 & ~n5304;
  assign n5406 = ~n1484 & ~n2706;
  assign n5407 = n5405 & n5406;
  assign n5408 = n5404 & n5407;
  assign n5409 = n5012 & n5408;
  assign n5410 = n457 & n5409;
  assign n5411 = n5392 & n5410;
  assign n5412 = n5381 & n5411;
  assign n5413 = n1122 & n5412;
  assign po79 = ~n5373 | ~n5413;
  assign n5415 = ~n590 & ~n2220;
  assign n5416 = ~pi020 & n5353;
  assign n5417 = n1044 & n1882;
  assign n5418 = ~n1697 & ~n5417;
  assign n5419 = ~n5416 & n5418;
  assign n5420 = n3677 & n5419;
  assign n5421 = n5415 & n5420;
  assign n5422 = n278 & n5397;
  assign n5423 = ~pi003 & ~n3502;
  assign n5424 = n1093 & ~n5423;
  assign n5425 = ~n5422 & n5424;
  assign n5426 = n1201 & n2200;
  assign n5427 = ~n1190 & ~n5426;
  assign n5428 = n3295 & n5427;
  assign n5429 = n5425 & n5428;
  assign n5430 = n5421 & n5429;
  assign n5431 = n5014 & n5430;
  assign n5432 = pi022 & n1694;
  assign n5433 = n466 & ~n5432;
  assign n5434 = ~n2036 & n3968;
  assign n5435 = n5433 & n5434;
  assign n5436 = n5431 & n5435;
  assign n5437 = ~n663 & ~n844;
  assign n5438 = n2227 & ~n5437;
  assign n5439 = n3867 & ~n5438;
  assign n5440 = n1558 & n5439;
  assign n5441 = n2991 & n5440;
  assign n5442 = n5436 & n5441;
  assign n5443 = n1660 & n5360;
  assign n5444 = ~n1797 & n5443;
  assign n5445 = n948 & n1414;
  assign n5446 = n494 & n1630;
  assign n5447 = n346 & n5446;
  assign n5448 = n3872 & ~n5447;
  assign n5449 = ~n5445 & n5448;
  assign n5450 = ~n1531 & ~n1676;
  assign n5451 = pi021 & ~n5450;
  assign n5452 = n1139 & ~n5451;
  assign n5453 = n3432 & n5452;
  assign n5454 = n5449 & n5453;
  assign n5455 = ~n383 & ~n5454;
  assign n5456 = n5444 & ~n5455;
  assign n5457 = n5349 & n5456;
  assign n5458 = n5371 & n5457;
  assign po80 = ~n5442 | ~n5458;
  assign n5460 = n1468 & ~n3041;
  assign n5461 = n1252 & ~n2124;
  assign n5462 = ~n2542 & n5461;
  assign n5463 = n5460 & n5462;
  assign n5464 = n1683 & n5463;
  assign n5465 = n1635 & n5307;
  assign n5466 = n5464 & n5465;
  assign n5467 = ~n1310 & n5444;
  assign n5468 = n5017 & n5467;
  assign n5469 = n1163 & n5468;
  assign n5470 = n2038 & n5469;
  assign po81 = ~n5466 | ~n5470;
  assign n5472 = ~n314 & ~n1018;
  assign n5473 = n4970 & n5472;
  assign n5474 = ~n298 & ~n331;
  assign n5475 = n1214 & n5474;
  assign n5476 = n3660 & n5475;
  assign n5477 = n1181 & n5476;
  assign po82 = ~n5473 | ~n5477;
  assign n5479 = ~n1471 & n3184;
  assign n5480 = ~n427 & n5479;
  assign n5481 = ~n323 & n5480;
  assign po83 = ~n1351 | ~n5481;
  assign po84 = ~n1322 | n1636;
  assign n5484 = n1433 & ~n4744;
  assign n5485 = ~n1070 & ~n5484;
  assign n5486 = ~n3803 & ~n4971;
  assign n5487 = ~po65 & n5486;
  assign po85 = n5485 | ~n5487;
  assign n5489 = n978 & n2291;
  assign n5490 = n2932 & ~n5489;
  assign n5491 = n230 & n4043;
  assign n5492 = ~n1476 & ~n5491;
  assign n5493 = ~n1521 & n5492;
  assign n5494 = n3602 & n5493;
  assign n5495 = ~n830 & n5494;
  assign n5496 = n5490 & n5495;
  assign po86 = ~n3495 | ~n5496;
  assign po87 = ~n4921 | po66;
  assign n5499 = pi023 & n2388;
  assign n5500 = ~n515 & n2886;
  assign n5501 = ~n5499 & ~n5500;
  assign n5502 = ~n2491 & ~n2492;
  assign n5503 = ~n2389 & n5502;
  assign n5504 = n4694 & n5503;
  assign n5505 = n1478 & n2333;
  assign n5506 = ~n1905 & ~n5505;
  assign n5507 = n2904 & n5506;
  assign n5508 = n5504 & n5507;
  assign n5509 = n5501 & n5508;
  assign n5510 = n3012 & ~n5489;
  assign n5511 = ~n2400 & ~n2948;
  assign n5512 = pi015 & ~n5511;
  assign n5513 = ~n2634 & ~n5512;
  assign n5514 = n5510 & n5513;
  assign n5515 = n3662 & n5514;
  assign n5516 = n5044 & n5515;
  assign n5517 = n5509 & n5516;
  assign po88 = ~n2443 | ~n5517;
  assign n5519 = n632 & n855;
  assign n5520 = pi019 & n1134;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = ~n4791 & n5521;
  assign n5523 = n4866 & ~n5522;
  assign n5524 = n4901 & ~n5523;
  assign n5525 = n2679 & n5524;
  assign n5526 = n4897 & n5525;
  assign n5527 = ~n1182 & ~n4453;
  assign n5528 = n3184 & n5527;
  assign n5529 = ~n4200 & n5528;
  assign n5530 = ~n595 & ~n599;
  assign n5531 = ~n302 & ~n1032;
  assign n5532 = n5530 & ~n5531;
  assign n5533 = n5529 & n5532;
  assign n5534 = n4222 & n5533;
  assign n5535 = n991 & n5484;
  assign n5536 = n1059 & ~n5535;
  assign n5537 = n702 & n1208;
  assign n5538 = n1930 & n5537;
  assign n5539 = ~n5536 & ~n5538;
  assign n5540 = n5534 & n5539;
  assign n5541 = n5526 & n5540;
  assign po89 = ~n4885 | ~n5541;
  assign n5543 = n4679 & n5490;
  assign n5544 = ~n3659 & n5543;
  assign po90 = ~n2443 | ~n5544;
  assign po91 = ~n1027 | ~n4987;
  assign n5547 = ~pi108 & n2309;
  assign po93 = ~n2792 | n5547;
  assign po40 = po27;
  assign po74 = po73;
  assign po75 = po73;
  assign po76 = po73;
endmodule


